-- soc_system.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		clk_clk                               : in    std_logic                     := '0';             --                       clk.clk
		hps_0_f2h_cold_reset_req_reset_n      : in    std_logic                     := '0';             --  hps_0_f2h_cold_reset_req.reset_n
		hps_0_f2h_debug_reset_req_reset_n     : in    std_logic                     := '0';             -- hps_0_f2h_debug_reset_req.reset_n
		hps_0_f2h_stm_hw_events_stm_hwevents  : in    std_logic_vector(27 downto 0) := (others => '0'); --   hps_0_f2h_stm_hw_events.stm_hwevents
		hps_0_f2h_warm_reset_req_reset_n      : in    std_logic                     := '0';             --  hps_0_f2h_warm_reset_req.reset_n
		hps_0_h2f_reset_reset_n               : out   std_logic;                                        --           hps_0_h2f_reset.reset_n
		hps_0_hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        --              hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		hps_0_hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --                          .hps_io_emac1_inst_TXD0
		hps_0_hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --                          .hps_io_emac1_inst_TXD1
		hps_0_hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --                          .hps_io_emac1_inst_TXD2
		hps_0_hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --                          .hps_io_emac1_inst_TXD3
		hps_0_hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RXD0
		hps_0_hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --                          .hps_io_emac1_inst_MDIO
		hps_0_hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --                          .hps_io_emac1_inst_MDC
		hps_0_hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RX_CTL
		hps_0_hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --                          .hps_io_emac1_inst_TX_CTL
		hps_0_hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RX_CLK
		hps_0_hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RXD1
		hps_0_hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RXD2
		hps_0_hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RXD3
		hps_0_hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_CMD
		hps_0_hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_D0
		hps_0_hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_D1
		hps_0_hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --                          .hps_io_sdio_inst_CLK
		hps_0_hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_D2
		hps_0_hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D0      : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D0
		hps_0_hps_io_hps_io_usb1_inst_D1      : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D1
		hps_0_hps_io_hps_io_usb1_inst_D2      : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D2
		hps_0_hps_io_hps_io_usb1_inst_D3      : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D4      : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D4
		hps_0_hps_io_hps_io_usb1_inst_D5      : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D5
		hps_0_hps_io_hps_io_usb1_inst_D6      : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D6
		hps_0_hps_io_hps_io_usb1_inst_D7      : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D7
		hps_0_hps_io_hps_io_usb1_inst_CLK     : in    std_logic                     := '0';             --                          .hps_io_usb1_inst_CLK
		hps_0_hps_io_hps_io_usb1_inst_STP     : out   std_logic;                                        --                          .hps_io_usb1_inst_STP
		hps_0_hps_io_hps_io_usb1_inst_DIR     : in    std_logic                     := '0';             --                          .hps_io_usb1_inst_DIR
		hps_0_hps_io_hps_io_usb1_inst_NXT     : in    std_logic                     := '0';             --                          .hps_io_usb1_inst_NXT
		hps_0_hps_io_hps_io_spim1_inst_CLK    : out   std_logic;                                        --                          .hps_io_spim1_inst_CLK
		hps_0_hps_io_hps_io_spim1_inst_MOSI   : out   std_logic;                                        --                          .hps_io_spim1_inst_MOSI
		hps_0_hps_io_hps_io_spim1_inst_MISO   : in    std_logic                     := '0';             --                          .hps_io_spim1_inst_MISO
		hps_0_hps_io_hps_io_spim1_inst_SS0    : out   std_logic;                                        --                          .hps_io_spim1_inst_SS0
		hps_0_hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --                          .hps_io_uart0_inst_RX
		hps_0_hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --                          .hps_io_uart0_inst_TX
		hps_0_hps_io_hps_io_i2c0_inst_SDA     : inout std_logic                     := '0';             --                          .hps_io_i2c0_inst_SDA
		hps_0_hps_io_hps_io_i2c0_inst_SCL     : inout std_logic                     := '0';             --                          .hps_io_i2c0_inst_SCL
		hps_0_hps_io_hps_io_i2c1_inst_SDA     : inout std_logic                     := '0';             --                          .hps_io_i2c1_inst_SDA
		hps_0_hps_io_hps_io_i2c1_inst_SCL     : inout std_logic                     := '0';             --                          .hps_io_i2c1_inst_SCL
		hps_0_hps_io_hps_io_gpio_inst_GPIO09  : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO09
		hps_0_hps_io_hps_io_gpio_inst_GPIO35  : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO35
		hps_0_hps_io_hps_io_gpio_inst_GPIO40  : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO40
		hps_0_hps_io_hps_io_gpio_inst_GPIO53  : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO53
		hps_0_hps_io_hps_io_gpio_inst_GPIO54  : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO54
		hps_0_hps_io_hps_io_gpio_inst_GPIO61  : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO61
		memory_mem_a                          : out   std_logic_vector(14 downto 0);                    --                    memory.mem_a
		memory_mem_ba                         : out   std_logic_vector(2 downto 0);                     --                          .mem_ba
		memory_mem_ck                         : out   std_logic;                                        --                          .mem_ck
		memory_mem_ck_n                       : out   std_logic;                                        --                          .mem_ck_n
		memory_mem_cke                        : out   std_logic;                                        --                          .mem_cke
		memory_mem_cs_n                       : out   std_logic;                                        --                          .mem_cs_n
		memory_mem_ras_n                      : out   std_logic;                                        --                          .mem_ras_n
		memory_mem_cas_n                      : out   std_logic;                                        --                          .mem_cas_n
		memory_mem_we_n                       : out   std_logic;                                        --                          .mem_we_n
		memory_mem_reset_n                    : out   std_logic;                                        --                          .mem_reset_n
		memory_mem_dq                         : inout std_logic_vector(31 downto 0) := (others => '0'); --                          .mem_dq
		memory_mem_dqs                        : inout std_logic_vector(3 downto 0)  := (others => '0'); --                          .mem_dqs
		memory_mem_dqs_n                      : inout std_logic_vector(3 downto 0)  := (others => '0'); --                          .mem_dqs_n
		memory_mem_odt                        : out   std_logic;                                        --                          .mem_odt
		memory_mem_dm                         : out   std_logic_vector(3 downto 0);                     --                          .mem_dm
		memory_oct_rzqin                      : in    std_logic                     := '0';             --                          .oct_rzqin
		reset_reset_n                         : in    std_logic                     := '0'              --                     reset.reset_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component soc_system_KBandIPsub is
		port (
			clk_clk                  : in  std_logic                      := 'X';             -- clk
			clk_int_clk              : in  std_logic                      := 'X';             -- clk
			kbandinput_1_csr_irq_irq : out std_logic;                                         -- irq
			kbandinput_2_csr_irq_irq : out std_logic;                                         -- irq
			kbandoutput_csr_irq_irq  : out std_logic;                                         -- irq
			m0_waitrequest           : in  std_logic                      := 'X';             -- waitrequest
			m0_readdata              : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid         : in  std_logic                      := 'X';             -- readdatavalid
			m0_burstcount            : out std_logic_vector(4 downto 0);                      -- burstcount
			m0_writedata             : out std_logic_vector(127 downto 0);                    -- writedata
			m0_address               : out std_logic_vector(29 downto 0);                     -- address
			m0_write                 : out std_logic;                                         -- write
			m0_read                  : out std_logic;                                         -- read
			m0_byteenable            : out std_logic_vector(15 downto 0);                     -- byteenable
			m0_debugaccess           : out std_logic;                                         -- debugaccess
			reset_reset_n            : in  std_logic                      := 'X';             -- reset_n
			sfpga_waitrequest        : out std_logic;                                         -- waitrequest
			sfpga_readdata           : out std_logic_vector(63 downto 0);                     -- readdata
			sfpga_readdatavalid      : out std_logic;                                         -- readdatavalid
			sfpga_burstcount         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- burstcount
			sfpga_writedata          : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- writedata
			sfpga_address            : in  std_logic_vector(17 downto 0)  := (others => 'X'); -- address
			sfpga_write              : in  std_logic                      := 'X';             -- write
			sfpga_read               : in  std_logic                      := 'X';             -- read
			sfpga_byteenable         : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- byteenable
			sfpga_debugaccess        : in  std_logic                      := 'X';             -- debugaccess
			slw_waitrequest          : out std_logic;                                         -- waitrequest
			slw_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			slw_readdatavalid        : out std_logic;                                         -- readdatavalid
			slw_burstcount           : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- burstcount
			slw_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			slw_address              : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- address
			slw_write                : in  std_logic                      := 'X';             -- write
			slw_read                 : in  std_logic                      := 'X';             -- read
			slw_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			slw_debugaccess          : in  std_logic                      := 'X'              -- debugaccess
		);
	end component soc_system_KBandIPsub;

	component axi_bridge_for_acp_128 is
		port (
			clk            : in  std_logic                      := 'X';             -- clk
			reset          : in  std_logic                      := 'X';             -- reset
			axm_m0_araddr  : out std_logic_vector(31 downto 0);                     -- araddr
			axm_m0_arburst : out std_logic_vector(1 downto 0);                      -- arburst
			axm_m0_arcache : out std_logic_vector(3 downto 0);                      -- arcache
			axm_m0_arid    : out std_logic_vector(7 downto 0);                      -- arid
			axm_m0_arlen   : out std_logic_vector(3 downto 0);                      -- arlen
			axm_m0_arlock  : out std_logic_vector(1 downto 0);                      -- arlock
			axm_m0_arprot  : out std_logic_vector(2 downto 0);                      -- arprot
			axm_m0_arready : in  std_logic                      := 'X';             -- arready
			axm_m0_arsize  : out std_logic_vector(2 downto 0);                      -- arsize
			axm_m0_aruser  : out std_logic_vector(4 downto 0);                      -- aruser
			axm_m0_arvalid : out std_logic;                                         -- arvalid
			axm_m0_awaddr  : out std_logic_vector(31 downto 0);                     -- awaddr
			axm_m0_awburst : out std_logic_vector(1 downto 0);                      -- awburst
			axm_m0_awcache : out std_logic_vector(3 downto 0);                      -- awcache
			axm_m0_awid    : out std_logic_vector(7 downto 0);                      -- awid
			axm_m0_awlen   : out std_logic_vector(3 downto 0);                      -- awlen
			axm_m0_awlock  : out std_logic_vector(1 downto 0);                      -- awlock
			axm_m0_awprot  : out std_logic_vector(2 downto 0);                      -- awprot
			axm_m0_awready : in  std_logic                      := 'X';             -- awready
			axm_m0_awsize  : out std_logic_vector(2 downto 0);                      -- awsize
			axm_m0_awuser  : out std_logic_vector(4 downto 0);                      -- awuser
			axm_m0_awvalid : out std_logic;                                         -- awvalid
			axm_m0_bid     : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- bid
			axm_m0_bready  : out std_logic;                                         -- bready
			axm_m0_bresp   : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			axm_m0_bvalid  : in  std_logic                      := 'X';             -- bvalid
			axm_m0_rdata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			axm_m0_rid     : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rid
			axm_m0_rlast   : in  std_logic                      := 'X';             -- rlast
			axm_m0_rready  : out std_logic;                                         -- rready
			axm_m0_rresp   : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			axm_m0_rvalid  : in  std_logic                      := 'X';             -- rvalid
			axm_m0_wdata   : out std_logic_vector(127 downto 0);                    -- wdata
			axm_m0_wid     : out std_logic_vector(7 downto 0);                      -- wid
			axm_m0_wlast   : out std_logic;                                         -- wlast
			axm_m0_wready  : in  std_logic                      := 'X';             -- wready
			axm_m0_wstrb   : out std_logic_vector(15 downto 0);                     -- wstrb
			axm_m0_wvalid  : out std_logic;                                         -- wvalid
			axs_s0_araddr  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			axs_s0_arburst : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			axs_s0_arcache : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			axs_s0_arid    : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			axs_s0_arlen   : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			axs_s0_arlock  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			axs_s0_arprot  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			axs_s0_arready : out std_logic;                                         -- arready
			axs_s0_arsize  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			axs_s0_aruser  : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			axs_s0_arvalid : in  std_logic                      := 'X';             -- arvalid
			axs_s0_awaddr  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			axs_s0_awburst : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			axs_s0_awcache : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			axs_s0_awid    : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			axs_s0_awlen   : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			axs_s0_awlock  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			axs_s0_awprot  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			axs_s0_awready : out std_logic;                                         -- awready
			axs_s0_awsize  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			axs_s0_awuser  : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			axs_s0_awvalid : in  std_logic                      := 'X';             -- awvalid
			axs_s0_bid     : out std_logic_vector(7 downto 0);                      -- bid
			axs_s0_bready  : in  std_logic                      := 'X';             -- bready
			axs_s0_bresp   : out std_logic_vector(1 downto 0);                      -- bresp
			axs_s0_bvalid  : out std_logic;                                         -- bvalid
			axs_s0_rdata   : out std_logic_vector(127 downto 0);                    -- rdata
			axs_s0_rid     : out std_logic_vector(7 downto 0);                      -- rid
			axs_s0_rlast   : out std_logic;                                         -- rlast
			axs_s0_rready  : in  std_logic                      := 'X';             -- rready
			axs_s0_rresp   : out std_logic_vector(1 downto 0);                      -- rresp
			axs_s0_rvalid  : out std_logic;                                         -- rvalid
			axs_s0_wdata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			axs_s0_wid     : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			axs_s0_wlast   : in  std_logic                      := 'X';             -- wlast
			axs_s0_wready  : out std_logic;                                         -- wready
			axs_s0_wstrb   : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			axs_s0_wvalid  : in  std_logic                      := 'X'              -- wvalid
		);
	end component axi_bridge_for_acp_128;

	component altera_address_span_extender is
		generic (
			DATA_WIDTH           : integer                       := 32;
			BYTEENABLE_WIDTH     : integer                       := 4;
			MASTER_ADDRESS_WIDTH : integer                       := 32;
			SLAVE_ADDRESS_WIDTH  : integer                       := 16;
			SLAVE_ADDRESS_SHIFT  : integer                       := 2;
			BURSTCOUNT_WIDTH     : integer                       := 1;
			CNTL_ADDRESS_WIDTH   : integer                       := 1;
			SUB_WINDOW_COUNT     : integer                       := 1;
			MASTER_ADDRESS_DEF   : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000"
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			avs_s0_address       : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			avs_s0_read          : in  std_logic                      := 'X';             -- read
			avs_s0_readdata      : out std_logic_vector(127 downto 0);                    -- readdata
			avs_s0_write         : in  std_logic                      := 'X';             -- write
			avs_s0_writedata     : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			avs_s0_readdatavalid : out std_logic;                                         -- readdatavalid
			avs_s0_waitrequest   : out std_logic;                                         -- waitrequest
			avs_s0_byteenable    : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			avs_s0_burstcount    : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- burstcount
			avm_m0_address       : out std_logic_vector(31 downto 0);                     -- address
			avm_m0_read          : out std_logic;                                         -- read
			avm_m0_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			avm_m0_readdata      : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			avm_m0_write         : out std_logic;                                         -- write
			avm_m0_writedata     : out std_logic_vector(127 downto 0);                    -- writedata
			avm_m0_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			avm_m0_byteenable    : out std_logic_vector(15 downto 0);                     -- byteenable
			avm_m0_burstcount    : out std_logic_vector(4 downto 0);                      -- burstcount
			avs_cntl_read        : in  std_logic                      := 'X';             -- read
			avs_cntl_readdata    : out std_logic_vector(63 downto 0);                     -- readdata
			avs_cntl_write       : in  std_logic                      := 'X';             -- write
			avs_cntl_writedata   : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- writedata
			avs_cntl_byteenable  : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- byteenable
			avs_cntl_address     : in  std_logic_vector(0 downto 0)   := (others => 'X')  -- address
		);
	end component altera_address_span_extender;

	component soc_system_fpga_only_master is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component soc_system_fpga_only_master;

	component soc_system_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			f2h_cold_rst_req_n       : in    std_logic                      := 'X';             -- reset_n
			f2h_dbg_rst_req_n        : in    std_logic                      := 'X';             -- reset_n
			f2h_warm_rst_req_n       : in    std_logic                      := 'X';             -- reset_n
			h2f_user0_clk            : out   std_logic;                                         -- clk
			h2f_user1_clk            : out   std_logic;                                         -- clk
			f2h_stm_hwevents         : in    std_logic_vector(27 downto 0)  := (others => 'X'); -- stm_hwevents
			mem_a                    : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                   : out   std_logic;                                         -- mem_ck
			mem_ck_n                 : out   std_logic;                                         -- mem_ck_n
			mem_cke                  : out   std_logic;                                         -- mem_cke
			mem_cs_n                 : out   std_logic;                                         -- mem_cs_n
			mem_ras_n                : out   std_logic;                                         -- mem_ras_n
			mem_cas_n                : out   std_logic;                                         -- mem_cas_n
			mem_we_n                 : out   std_logic;                                         -- mem_we_n
			mem_reset_n              : out   std_logic;                                         -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                         -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin                : in    std_logic                      := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                         -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                         -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                         -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                         -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                         -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                      := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                         -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                         -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                      := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                         -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                         -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                         -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                         -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                      := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                         -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                      := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                         -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                         -- reset_n
			f2h_sdram0_clk           : in    std_logic                      := 'X';             -- clk
			f2h_sdram0_ADDRESS       : in    std_logic_vector(26 downto 0)  := (others => 'X'); -- address
			f2h_sdram0_BURSTCOUNT    : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			f2h_sdram0_WAITREQUEST   : out   std_logic;                                         -- waitrequest
			f2h_sdram0_READDATA      : out   std_logic_vector(255 downto 0);                    -- readdata
			f2h_sdram0_READDATAVALID : out   std_logic;                                         -- readdatavalid
			f2h_sdram0_READ          : in    std_logic                      := 'X';             -- read
			f2h_sdram0_WRITEDATA     : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			f2h_sdram0_BYTEENABLE    : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			f2h_sdram0_WRITE         : in    std_logic                      := 'X';             -- write
			h2f_axi_clk              : in    std_logic                      := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID              : out   std_logic;                                         -- awvalid
			h2f_AWREADY              : in    std_logic                      := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA                : out   std_logic_vector(63 downto 0);                     -- wdata
			h2f_WSTRB                : out   std_logic_vector(7 downto 0);                      -- wstrb
			h2f_WLAST                : out   std_logic;                                         -- wlast
			h2f_WVALID               : out   std_logic;                                         -- wvalid
			h2f_WREADY               : in    std_logic                      := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                         -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID              : out   std_logic;                                         -- arvalid
			h2f_ARREADY              : in    std_logic                      := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(63 downto 0)  := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                         -- rready
			f2h_axi_clk              : in    std_logic                      := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                         -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                         -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID               : out   std_logic;                                         -- bvalid
			f2h_BREADY               : in    std_logic                      := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                         -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA                : out   std_logic_vector(127 downto 0);                    -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST                : out   std_logic;                                         -- rlast
			f2h_RVALID               : out   std_logic;                                         -- rvalid
			f2h_RREADY               : in    std_logic                      := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY           : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                         -- wlast
			h2f_lw_WVALID            : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY            : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                         -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY           : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                         -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0)  := (others => 'X')  -- irq
		);
	end component soc_system_hps_0;

	component intr_capturer is
		generic (
			NUM_INTR : integer := 32
		);
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			rst_n        : in  std_logic                     := 'X';             -- reset_n
			addr         : in  std_logic                     := 'X';             -- address
			read         : in  std_logic                     := 'X';             -- read
			rddata       : out std_logic_vector(31 downto 0);                    -- readdata
			interrupt_in : in  std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component intr_capturer;

	component soc_system_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component soc_system_pll_0;

	component soc_system_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_sysid_qsys;

	component soc_system_mm_interconnect_0 is
		port (
			axi_bridge_for_acp_128_0_s0_awid                 : out std_logic_vector(7 downto 0);                      -- awid
			axi_bridge_for_acp_128_0_s0_awaddr               : out std_logic_vector(31 downto 0);                     -- awaddr
			axi_bridge_for_acp_128_0_s0_awlen                : out std_logic_vector(3 downto 0);                      -- awlen
			axi_bridge_for_acp_128_0_s0_awsize               : out std_logic_vector(2 downto 0);                      -- awsize
			axi_bridge_for_acp_128_0_s0_awburst              : out std_logic_vector(1 downto 0);                      -- awburst
			axi_bridge_for_acp_128_0_s0_awlock               : out std_logic_vector(1 downto 0);                      -- awlock
			axi_bridge_for_acp_128_0_s0_awcache              : out std_logic_vector(3 downto 0);                      -- awcache
			axi_bridge_for_acp_128_0_s0_awprot               : out std_logic_vector(2 downto 0);                      -- awprot
			axi_bridge_for_acp_128_0_s0_awuser               : out std_logic_vector(4 downto 0);                      -- awuser
			axi_bridge_for_acp_128_0_s0_awvalid              : out std_logic;                                         -- awvalid
			axi_bridge_for_acp_128_0_s0_awready              : in  std_logic                      := 'X';             -- awready
			axi_bridge_for_acp_128_0_s0_wid                  : out std_logic_vector(7 downto 0);                      -- wid
			axi_bridge_for_acp_128_0_s0_wdata                : out std_logic_vector(127 downto 0);                    -- wdata
			axi_bridge_for_acp_128_0_s0_wstrb                : out std_logic_vector(15 downto 0);                     -- wstrb
			axi_bridge_for_acp_128_0_s0_wlast                : out std_logic;                                         -- wlast
			axi_bridge_for_acp_128_0_s0_wvalid               : out std_logic;                                         -- wvalid
			axi_bridge_for_acp_128_0_s0_wready               : in  std_logic                      := 'X';             -- wready
			axi_bridge_for_acp_128_0_s0_bid                  : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- bid
			axi_bridge_for_acp_128_0_s0_bresp                : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			axi_bridge_for_acp_128_0_s0_bvalid               : in  std_logic                      := 'X';             -- bvalid
			axi_bridge_for_acp_128_0_s0_bready               : out std_logic;                                         -- bready
			axi_bridge_for_acp_128_0_s0_arid                 : out std_logic_vector(7 downto 0);                      -- arid
			axi_bridge_for_acp_128_0_s0_araddr               : out std_logic_vector(31 downto 0);                     -- araddr
			axi_bridge_for_acp_128_0_s0_arlen                : out std_logic_vector(3 downto 0);                      -- arlen
			axi_bridge_for_acp_128_0_s0_arsize               : out std_logic_vector(2 downto 0);                      -- arsize
			axi_bridge_for_acp_128_0_s0_arburst              : out std_logic_vector(1 downto 0);                      -- arburst
			axi_bridge_for_acp_128_0_s0_arlock               : out std_logic_vector(1 downto 0);                      -- arlock
			axi_bridge_for_acp_128_0_s0_arcache              : out std_logic_vector(3 downto 0);                      -- arcache
			axi_bridge_for_acp_128_0_s0_arprot               : out std_logic_vector(2 downto 0);                      -- arprot
			axi_bridge_for_acp_128_0_s0_aruser               : out std_logic_vector(4 downto 0);                      -- aruser
			axi_bridge_for_acp_128_0_s0_arvalid              : out std_logic;                                         -- arvalid
			axi_bridge_for_acp_128_0_s0_arready              : in  std_logic                      := 'X';             -- arready
			axi_bridge_for_acp_128_0_s0_rid                  : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rid
			axi_bridge_for_acp_128_0_s0_rdata                : in  std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			axi_bridge_for_acp_128_0_s0_rresp                : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			axi_bridge_for_acp_128_0_s0_rlast                : in  std_logic                      := 'X';             -- rlast
			axi_bridge_for_acp_128_0_s0_rvalid               : in  std_logic                      := 'X';             -- rvalid
			axi_bridge_for_acp_128_0_s0_rready               : out std_logic;                                         -- rready
			pll_0_outclk0_clk                                : in  std_logic                      := 'X';             -- clk
			fft_ddr_bridge_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			fft_ddr_bridge_expanded_master_address           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			fft_ddr_bridge_expanded_master_waitrequest       : out std_logic;                                         -- waitrequest
			fft_ddr_bridge_expanded_master_burstcount        : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- burstcount
			fft_ddr_bridge_expanded_master_byteenable        : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			fft_ddr_bridge_expanded_master_read              : in  std_logic                      := 'X';             -- read
			fft_ddr_bridge_expanded_master_readdata          : out std_logic_vector(127 downto 0);                    -- readdata
			fft_ddr_bridge_expanded_master_readdatavalid     : out std_logic;                                         -- readdatavalid
			fft_ddr_bridge_expanded_master_write             : in  std_logic                      := 'X';             -- write
			fft_ddr_bridge_expanded_master_writedata         : in  std_logic_vector(127 downto 0) := (others => 'X')  -- writedata
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_mm_interconnect_1 is
		port (
			hps_0_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_axi_master_wdata                                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_axi_master_wstrb                                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_axi_master_rdata                                       : out std_logic_vector(63 downto 0);                    -- rdata
			hps_0_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			pll_0_outclk0_clk                                                : in  std_logic                     := 'X';             -- clk
			FPGA_Slave_mm_bridge_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			FPGA_Slave_mm_bridge_s0_address                                  : out std_logic_vector(17 downto 0);                    -- address
			FPGA_Slave_mm_bridge_s0_write                                    : out std_logic;                                        -- write
			FPGA_Slave_mm_bridge_s0_read                                     : out std_logic;                                        -- read
			FPGA_Slave_mm_bridge_s0_readdata                                 : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			FPGA_Slave_mm_bridge_s0_writedata                                : out std_logic_vector(63 downto 0);                    -- writedata
			FPGA_Slave_mm_bridge_s0_burstcount                               : out std_logic_vector(0 downto 0);                     -- burstcount
			FPGA_Slave_mm_bridge_s0_byteenable                               : out std_logic_vector(7 downto 0);                     -- byteenable
			FPGA_Slave_mm_bridge_s0_readdatavalid                            : in  std_logic                     := 'X';             -- readdatavalid
			FPGA_Slave_mm_bridge_s0_waitrequest                              : in  std_logic                     := 'X';             -- waitrequest
			FPGA_Slave_mm_bridge_s0_debugaccess                              : out std_logic                                         -- debugaccess
		);
	end component soc_system_mm_interconnect_1;

	component soc_system_mm_interconnect_2 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			pll_0_outclk0_clk                                                   : in  std_logic                     := 'X';             -- clk
			fpga_only_master_clk_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			lw_mm_bridge_reset_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			fpga_only_master_master_address                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			fpga_only_master_master_waitrequest                                 : out std_logic;                                        -- waitrequest
			fpga_only_master_master_byteenable                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			fpga_only_master_master_read                                        : in  std_logic                     := 'X';             -- read
			fpga_only_master_master_readdata                                    : out std_logic_vector(31 downto 0);                    -- readdata
			fpga_only_master_master_readdatavalid                               : out std_logic;                                        -- readdatavalid
			fpga_only_master_master_write                                       : in  std_logic                     := 'X';             -- write
			fpga_only_master_master_writedata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			lw_mm_bridge_s0_address                                             : out std_logic_vector(19 downto 0);                    -- address
			lw_mm_bridge_s0_write                                               : out std_logic;                                        -- write
			lw_mm_bridge_s0_read                                                : out std_logic;                                        -- read
			lw_mm_bridge_s0_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			lw_mm_bridge_s0_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			lw_mm_bridge_s0_burstcount                                          : out std_logic_vector(0 downto 0);                     -- burstcount
			lw_mm_bridge_s0_byteenable                                          : out std_logic_vector(3 downto 0);                     -- byteenable
			lw_mm_bridge_s0_readdatavalid                                       : in  std_logic                     := 'X';             -- readdatavalid
			lw_mm_bridge_s0_waitrequest                                         : in  std_logic                     := 'X';             -- waitrequest
			lw_mm_bridge_s0_debugaccess                                         : out std_logic                                         -- debugaccess
		);
	end component soc_system_mm_interconnect_2;

	component soc_system_mm_interconnect_3 is
		port (
			pll_0_outclk0_clk                              : in  std_logic                     := 'X';             -- clk
			KBandIPsub_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			lw_mm_bridge_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			lw_mm_bridge_m0_address                        : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			lw_mm_bridge_m0_waitrequest                    : out std_logic;                                        -- waitrequest
			lw_mm_bridge_m0_burstcount                     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			lw_mm_bridge_m0_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			lw_mm_bridge_m0_read                           : in  std_logic                     := 'X';             -- read
			lw_mm_bridge_m0_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			lw_mm_bridge_m0_readdatavalid                  : out std_logic;                                        -- readdatavalid
			lw_mm_bridge_m0_write                          : in  std_logic                     := 'X';             -- write
			lw_mm_bridge_m0_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			lw_mm_bridge_m0_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			intr_capturer_0_avalon_slave_0_address         : out std_logic_vector(0 downto 0);                     -- address
			intr_capturer_0_avalon_slave_0_read            : out std_logic;                                        -- read
			intr_capturer_0_avalon_slave_0_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			KBandIPsub_slw_address                         : out std_logic_vector(16 downto 0);                    -- address
			KBandIPsub_slw_write                           : out std_logic;                                        -- write
			KBandIPsub_slw_read                            : out std_logic;                                        -- read
			KBandIPsub_slw_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			KBandIPsub_slw_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			KBandIPsub_slw_burstcount                      : out std_logic_vector(0 downto 0);                     -- burstcount
			KBandIPsub_slw_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			KBandIPsub_slw_readdatavalid                   : in  std_logic                     := 'X';             -- readdatavalid
			KBandIPsub_slw_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			KBandIPsub_slw_debugaccess                     : out std_logic;                                        -- debugaccess
			sysid_qsys_control_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_mm_interconnect_3;

	component soc_system_mm_interconnect_6 is
		port (
			pll_0_outclk0_clk                                : in  std_logic                      := 'X';             -- clk
			fft_ddr_bridge_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			KBandIPsub_reset_reset_bridge_in_reset_reset     : in  std_logic                      := 'X';             -- reset
			KBandIPsub_m0_address                            : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- address
			KBandIPsub_m0_waitrequest                        : out std_logic;                                         -- waitrequest
			KBandIPsub_m0_burstcount                         : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- burstcount
			KBandIPsub_m0_byteenable                         : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			KBandIPsub_m0_read                               : in  std_logic                      := 'X';             -- read
			KBandIPsub_m0_readdata                           : out std_logic_vector(127 downto 0);                    -- readdata
			KBandIPsub_m0_readdatavalid                      : out std_logic;                                         -- readdatavalid
			KBandIPsub_m0_write                              : in  std_logic                      := 'X';             -- write
			KBandIPsub_m0_writedata                          : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			KBandIPsub_m0_debugaccess                        : in  std_logic                      := 'X';             -- debugaccess
			fft_ddr_bridge_windowed_slave_address            : out std_logic_vector(25 downto 0);                     -- address
			fft_ddr_bridge_windowed_slave_write              : out std_logic;                                         -- write
			fft_ddr_bridge_windowed_slave_read               : out std_logic;                                         -- read
			fft_ddr_bridge_windowed_slave_readdata           : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			fft_ddr_bridge_windowed_slave_writedata          : out std_logic_vector(127 downto 0);                    -- writedata
			fft_ddr_bridge_windowed_slave_burstcount         : out std_logic_vector(4 downto 0);                      -- burstcount
			fft_ddr_bridge_windowed_slave_byteenable         : out std_logic_vector(15 downto 0);                     -- byteenable
			fft_ddr_bridge_windowed_slave_readdatavalid      : in  std_logic                      := 'X';             -- readdatavalid
			fft_ddr_bridge_windowed_slave_waitrequest        : in  std_logic                      := 'X'              -- waitrequest
		);
	end component soc_system_mm_interconnect_6;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component soc_system_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper_001;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	component soc_system_fpga_slave_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(63 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(63 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(17 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(7 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component soc_system_fpga_slave_mm_bridge;

	component soc_system_lw_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(19 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component soc_system_lw_mm_bridge;

	signal axi_bridge_for_acp_128_0_m0_awburst                           : std_logic_vector(1 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_awburst -> hps_0:f2h_AWBURST
	signal axi_bridge_for_acp_128_0_m0_arlen                             : std_logic_vector(3 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_arlen -> hps_0:f2h_ARLEN
	signal axi_bridge_for_acp_128_0_m0_awuser                            : std_logic_vector(4 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_awuser -> hps_0:f2h_AWUSER
	signal axi_bridge_for_acp_128_0_m0_wready                            : std_logic;                      -- hps_0:f2h_WREADY -> axi_bridge_for_acp_128_0:axm_m0_wready
	signal axi_bridge_for_acp_128_0_m0_wstrb                             : std_logic_vector(15 downto 0);  -- axi_bridge_for_acp_128_0:axm_m0_wstrb -> hps_0:f2h_WSTRB
	signal axi_bridge_for_acp_128_0_m0_rid                               : std_logic_vector(7 downto 0);   -- hps_0:f2h_RID -> axi_bridge_for_acp_128_0:axm_m0_rid
	signal axi_bridge_for_acp_128_0_m0_rready                            : std_logic;                      -- axi_bridge_for_acp_128_0:axm_m0_rready -> hps_0:f2h_RREADY
	signal axi_bridge_for_acp_128_0_m0_awlen                             : std_logic_vector(3 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_awlen -> hps_0:f2h_AWLEN
	signal axi_bridge_for_acp_128_0_m0_wid                               : std_logic_vector(7 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_wid -> hps_0:f2h_WID
	signal axi_bridge_for_acp_128_0_m0_arcache                           : std_logic_vector(3 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_arcache -> hps_0:f2h_ARCACHE
	signal axi_bridge_for_acp_128_0_m0_araddr                            : std_logic_vector(31 downto 0);  -- axi_bridge_for_acp_128_0:axm_m0_araddr -> hps_0:f2h_ARADDR
	signal axi_bridge_for_acp_128_0_m0_wvalid                            : std_logic;                      -- axi_bridge_for_acp_128_0:axm_m0_wvalid -> hps_0:f2h_WVALID
	signal axi_bridge_for_acp_128_0_m0_arprot                            : std_logic_vector(2 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_arprot -> hps_0:f2h_ARPROT
	signal axi_bridge_for_acp_128_0_m0_arvalid                           : std_logic;                      -- axi_bridge_for_acp_128_0:axm_m0_arvalid -> hps_0:f2h_ARVALID
	signal axi_bridge_for_acp_128_0_m0_awprot                            : std_logic_vector(2 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_awprot -> hps_0:f2h_AWPROT
	signal axi_bridge_for_acp_128_0_m0_wdata                             : std_logic_vector(127 downto 0); -- axi_bridge_for_acp_128_0:axm_m0_wdata -> hps_0:f2h_WDATA
	signal axi_bridge_for_acp_128_0_m0_arid                              : std_logic_vector(7 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_arid -> hps_0:f2h_ARID
	signal axi_bridge_for_acp_128_0_m0_awcache                           : std_logic_vector(3 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_awcache -> hps_0:f2h_AWCACHE
	signal axi_bridge_for_acp_128_0_m0_arlock                            : std_logic_vector(1 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_arlock -> hps_0:f2h_ARLOCK
	signal axi_bridge_for_acp_128_0_m0_awlock                            : std_logic_vector(1 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_awlock -> hps_0:f2h_AWLOCK
	signal axi_bridge_for_acp_128_0_m0_awaddr                            : std_logic_vector(31 downto 0);  -- axi_bridge_for_acp_128_0:axm_m0_awaddr -> hps_0:f2h_AWADDR
	signal axi_bridge_for_acp_128_0_m0_arready                           : std_logic;                      -- hps_0:f2h_ARREADY -> axi_bridge_for_acp_128_0:axm_m0_arready
	signal axi_bridge_for_acp_128_0_m0_bresp                             : std_logic_vector(1 downto 0);   -- hps_0:f2h_BRESP -> axi_bridge_for_acp_128_0:axm_m0_bresp
	signal axi_bridge_for_acp_128_0_m0_rdata                             : std_logic_vector(127 downto 0); -- hps_0:f2h_RDATA -> axi_bridge_for_acp_128_0:axm_m0_rdata
	signal axi_bridge_for_acp_128_0_m0_arburst                           : std_logic_vector(1 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_arburst -> hps_0:f2h_ARBURST
	signal axi_bridge_for_acp_128_0_m0_awready                           : std_logic;                      -- hps_0:f2h_AWREADY -> axi_bridge_for_acp_128_0:axm_m0_awready
	signal axi_bridge_for_acp_128_0_m0_arsize                            : std_logic_vector(2 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_arsize -> hps_0:f2h_ARSIZE
	signal axi_bridge_for_acp_128_0_m0_bready                            : std_logic;                      -- axi_bridge_for_acp_128_0:axm_m0_bready -> hps_0:f2h_BREADY
	signal axi_bridge_for_acp_128_0_m0_rlast                             : std_logic;                      -- hps_0:f2h_RLAST -> axi_bridge_for_acp_128_0:axm_m0_rlast
	signal axi_bridge_for_acp_128_0_m0_wlast                             : std_logic;                      -- axi_bridge_for_acp_128_0:axm_m0_wlast -> hps_0:f2h_WLAST
	signal axi_bridge_for_acp_128_0_m0_rresp                             : std_logic_vector(1 downto 0);   -- hps_0:f2h_RRESP -> axi_bridge_for_acp_128_0:axm_m0_rresp
	signal axi_bridge_for_acp_128_0_m0_awid                              : std_logic_vector(7 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_awid -> hps_0:f2h_AWID
	signal axi_bridge_for_acp_128_0_m0_bid                               : std_logic_vector(7 downto 0);   -- hps_0:f2h_BID -> axi_bridge_for_acp_128_0:axm_m0_bid
	signal axi_bridge_for_acp_128_0_m0_bvalid                            : std_logic;                      -- hps_0:f2h_BVALID -> axi_bridge_for_acp_128_0:axm_m0_bvalid
	signal axi_bridge_for_acp_128_0_m0_aruser                            : std_logic_vector(4 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_aruser -> hps_0:f2h_ARUSER
	signal axi_bridge_for_acp_128_0_m0_awsize                            : std_logic_vector(2 downto 0);   -- axi_bridge_for_acp_128_0:axm_m0_awsize -> hps_0:f2h_AWSIZE
	signal axi_bridge_for_acp_128_0_m0_awvalid                           : std_logic;                      -- axi_bridge_for_acp_128_0:axm_m0_awvalid -> hps_0:f2h_AWVALID
	signal axi_bridge_for_acp_128_0_m0_rvalid                            : std_logic;                      -- hps_0:f2h_RVALID -> axi_bridge_for_acp_128_0:axm_m0_rvalid
	signal fpga_slave_mm_bridge_m0_waitrequest                           : std_logic;                      -- KBandIPsub:sfpga_waitrequest -> FPGA_Slave_mm_bridge:m0_waitrequest
	signal fpga_slave_mm_bridge_m0_readdata                              : std_logic_vector(63 downto 0);  -- KBandIPsub:sfpga_readdata -> FPGA_Slave_mm_bridge:m0_readdata
	signal fpga_slave_mm_bridge_m0_debugaccess                           : std_logic;                      -- FPGA_Slave_mm_bridge:m0_debugaccess -> KBandIPsub:sfpga_debugaccess
	signal fpga_slave_mm_bridge_m0_address                               : std_logic_vector(17 downto 0);  -- FPGA_Slave_mm_bridge:m0_address -> KBandIPsub:sfpga_address
	signal fpga_slave_mm_bridge_m0_read                                  : std_logic;                      -- FPGA_Slave_mm_bridge:m0_read -> KBandIPsub:sfpga_read
	signal fpga_slave_mm_bridge_m0_byteenable                            : std_logic_vector(7 downto 0);   -- FPGA_Slave_mm_bridge:m0_byteenable -> KBandIPsub:sfpga_byteenable
	signal fpga_slave_mm_bridge_m0_readdatavalid                         : std_logic;                      -- KBandIPsub:sfpga_readdatavalid -> FPGA_Slave_mm_bridge:m0_readdatavalid
	signal fpga_slave_mm_bridge_m0_writedata                             : std_logic_vector(63 downto 0);  -- FPGA_Slave_mm_bridge:m0_writedata -> KBandIPsub:sfpga_writedata
	signal fpga_slave_mm_bridge_m0_write                                 : std_logic;                      -- FPGA_Slave_mm_bridge:m0_write -> KBandIPsub:sfpga_write
	signal fpga_slave_mm_bridge_m0_burstcount                            : std_logic_vector(0 downto 0);   -- FPGA_Slave_mm_bridge:m0_burstcount -> KBandIPsub:sfpga_burstcount
	signal pll_0_outclk0_clk                                             : std_logic;                      -- pll_0:outclk_0 -> [FPGA_Slave_mm_bridge:clk, KBandIPsub:clk_clk, axi_bridge_for_acp_128_0:clk, fft_ddr_bridge:clk, fpga_only_master:clk_clk, hps_0:f2h_axi_clk, hps_0:f2h_sdram0_clk, hps_0:h2f_axi_clk, hps_0:h2f_lw_axi_clk, intr_capturer_0:clk, irq_mapper_002:clk, lw_mm_bridge:clk, mm_interconnect_0:pll_0_outclk0_clk, mm_interconnect_1:pll_0_outclk0_clk, mm_interconnect_2:pll_0_outclk0_clk, mm_interconnect_3:pll_0_outclk0_clk, mm_interconnect_6:pll_0_outclk0_clk, rst_controller:clk, rst_controller_001:clk, sysid_qsys:clock]
	signal pll_0_outclk1_clk                                             : std_logic;                      -- pll_0:outclk_1 -> KBandIPsub:clk_int_clk
	signal hps_0_h2f_reset_reset                                         : std_logic;                      -- hps_0:h2f_rst_n -> [hps_0_h2f_reset_reset_n, hps_0_h2f_reset_reset_n:in]
	signal fft_ddr_bridge_expanded_master_waitrequest                    : std_logic;                      -- mm_interconnect_0:fft_ddr_bridge_expanded_master_waitrequest -> fft_ddr_bridge:avm_m0_waitrequest
	signal fft_ddr_bridge_expanded_master_readdata                       : std_logic_vector(127 downto 0); -- mm_interconnect_0:fft_ddr_bridge_expanded_master_readdata -> fft_ddr_bridge:avm_m0_readdata
	signal fft_ddr_bridge_expanded_master_address                        : std_logic_vector(31 downto 0);  -- fft_ddr_bridge:avm_m0_address -> mm_interconnect_0:fft_ddr_bridge_expanded_master_address
	signal fft_ddr_bridge_expanded_master_read                           : std_logic;                      -- fft_ddr_bridge:avm_m0_read -> mm_interconnect_0:fft_ddr_bridge_expanded_master_read
	signal fft_ddr_bridge_expanded_master_byteenable                     : std_logic_vector(15 downto 0);  -- fft_ddr_bridge:avm_m0_byteenable -> mm_interconnect_0:fft_ddr_bridge_expanded_master_byteenable
	signal fft_ddr_bridge_expanded_master_readdatavalid                  : std_logic;                      -- mm_interconnect_0:fft_ddr_bridge_expanded_master_readdatavalid -> fft_ddr_bridge:avm_m0_readdatavalid
	signal fft_ddr_bridge_expanded_master_write                          : std_logic;                      -- fft_ddr_bridge:avm_m0_write -> mm_interconnect_0:fft_ddr_bridge_expanded_master_write
	signal fft_ddr_bridge_expanded_master_writedata                      : std_logic_vector(127 downto 0); -- fft_ddr_bridge:avm_m0_writedata -> mm_interconnect_0:fft_ddr_bridge_expanded_master_writedata
	signal fft_ddr_bridge_expanded_master_burstcount                     : std_logic_vector(4 downto 0);   -- fft_ddr_bridge:avm_m0_burstcount -> mm_interconnect_0:fft_ddr_bridge_expanded_master_burstcount
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awburst         : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awburst -> axi_bridge_for_acp_128_0:axs_s0_awburst
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awuser          : std_logic_vector(4 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awuser -> axi_bridge_for_acp_128_0:axs_s0_awuser
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlen           : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arlen -> axi_bridge_for_acp_128_0:axs_s0_arlen
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wstrb           : std_logic_vector(15 downto 0);  -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wstrb -> axi_bridge_for_acp_128_0:axs_s0_wstrb
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wready          : std_logic;                      -- axi_bridge_for_acp_128_0:axs_s0_wready -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wready
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rid             : std_logic_vector(7 downto 0);   -- axi_bridge_for_acp_128_0:axs_s0_rid -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rready          : std_logic;                      -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rready -> axi_bridge_for_acp_128_0:axs_s0_rready
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlen           : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awlen -> axi_bridge_for_acp_128_0:axs_s0_awlen
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wid             : std_logic_vector(7 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wid -> axi_bridge_for_acp_128_0:axs_s0_wid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arcache         : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arcache -> axi_bridge_for_acp_128_0:axs_s0_arcache
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wvalid          : std_logic;                      -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wvalid -> axi_bridge_for_acp_128_0:axs_s0_wvalid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_araddr          : std_logic_vector(31 downto 0);  -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_araddr -> axi_bridge_for_acp_128_0:axs_s0_araddr
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arprot          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arprot -> axi_bridge_for_acp_128_0:axs_s0_arprot
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awprot          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awprot -> axi_bridge_for_acp_128_0:axs_s0_awprot
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wdata           : std_logic_vector(127 downto 0); -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wdata -> axi_bridge_for_acp_128_0:axs_s0_wdata
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arvalid         : std_logic;                      -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arvalid -> axi_bridge_for_acp_128_0:axs_s0_arvalid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awcache         : std_logic_vector(3 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awcache -> axi_bridge_for_acp_128_0:axs_s0_awcache
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arid            : std_logic_vector(7 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arid -> axi_bridge_for_acp_128_0:axs_s0_arid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlock          : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arlock -> axi_bridge_for_acp_128_0:axs_s0_arlock
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlock          : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awlock -> axi_bridge_for_acp_128_0:axs_s0_awlock
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awaddr          : std_logic_vector(31 downto 0);  -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awaddr -> axi_bridge_for_acp_128_0:axs_s0_awaddr
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bresp           : std_logic_vector(1 downto 0);   -- axi_bridge_for_acp_128_0:axs_s0_bresp -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_bresp
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arready         : std_logic;                      -- axi_bridge_for_acp_128_0:axs_s0_arready -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arready
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rdata           : std_logic_vector(127 downto 0); -- axi_bridge_for_acp_128_0:axs_s0_rdata -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rdata
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awready         : std_logic;                      -- axi_bridge_for_acp_128_0:axs_s0_awready -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awready
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arburst         : std_logic_vector(1 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arburst -> axi_bridge_for_acp_128_0:axs_s0_arburst
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arsize          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arsize -> axi_bridge_for_acp_128_0:axs_s0_arsize
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bready          : std_logic;                      -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_bready -> axi_bridge_for_acp_128_0:axs_s0_bready
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rlast           : std_logic;                      -- axi_bridge_for_acp_128_0:axs_s0_rlast -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rlast
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wlast           : std_logic;                      -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wlast -> axi_bridge_for_acp_128_0:axs_s0_wlast
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rresp           : std_logic_vector(1 downto 0);   -- axi_bridge_for_acp_128_0:axs_s0_rresp -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rresp
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awid            : std_logic_vector(7 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awid -> axi_bridge_for_acp_128_0:axs_s0_awid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bid             : std_logic_vector(7 downto 0);   -- axi_bridge_for_acp_128_0:axs_s0_bid -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_bid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bvalid          : std_logic;                      -- axi_bridge_for_acp_128_0:axs_s0_bvalid -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_bvalid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awsize          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awsize -> axi_bridge_for_acp_128_0:axs_s0_awsize
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awvalid         : std_logic;                      -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awvalid -> axi_bridge_for_acp_128_0:axs_s0_awvalid
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_aruser          : std_logic_vector(4 downto 0);   -- mm_interconnect_0:axi_bridge_for_acp_128_0_s0_aruser -> axi_bridge_for_acp_128_0:axs_s0_aruser
	signal mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rvalid          : std_logic;                      -- axi_bridge_for_acp_128_0:axs_s0_rvalid -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rvalid
	signal hps_0_h2f_axi_master_awburst                                  : std_logic_vector(1 downto 0);   -- hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	signal hps_0_h2f_axi_master_arlen                                    : std_logic_vector(3 downto 0);   -- hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	signal hps_0_h2f_axi_master_wstrb                                    : std_logic_vector(7 downto 0);   -- hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	signal hps_0_h2f_axi_master_wready                                   : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	signal hps_0_h2f_axi_master_rid                                      : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	signal hps_0_h2f_axi_master_rready                                   : std_logic;                      -- hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	signal hps_0_h2f_axi_master_awlen                                    : std_logic_vector(3 downto 0);   -- hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	signal hps_0_h2f_axi_master_wid                                      : std_logic_vector(11 downto 0);  -- hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	signal hps_0_h2f_axi_master_arcache                                  : std_logic_vector(3 downto 0);   -- hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	signal hps_0_h2f_axi_master_wvalid                                   : std_logic;                      -- hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	signal hps_0_h2f_axi_master_araddr                                   : std_logic_vector(29 downto 0);  -- hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	signal hps_0_h2f_axi_master_arprot                                   : std_logic_vector(2 downto 0);   -- hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	signal hps_0_h2f_axi_master_awprot                                   : std_logic_vector(2 downto 0);   -- hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	signal hps_0_h2f_axi_master_wdata                                    : std_logic_vector(63 downto 0);  -- hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	signal hps_0_h2f_axi_master_arvalid                                  : std_logic;                      -- hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	signal hps_0_h2f_axi_master_awcache                                  : std_logic_vector(3 downto 0);   -- hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	signal hps_0_h2f_axi_master_arid                                     : std_logic_vector(11 downto 0);  -- hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	signal hps_0_h2f_axi_master_arlock                                   : std_logic_vector(1 downto 0);   -- hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	signal hps_0_h2f_axi_master_awlock                                   : std_logic_vector(1 downto 0);   -- hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	signal hps_0_h2f_axi_master_awaddr                                   : std_logic_vector(29 downto 0);  -- hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	signal hps_0_h2f_axi_master_bresp                                    : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	signal hps_0_h2f_axi_master_arready                                  : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	signal hps_0_h2f_axi_master_rdata                                    : std_logic_vector(63 downto 0);  -- mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	signal hps_0_h2f_axi_master_awready                                  : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	signal hps_0_h2f_axi_master_arburst                                  : std_logic_vector(1 downto 0);   -- hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	signal hps_0_h2f_axi_master_arsize                                   : std_logic_vector(2 downto 0);   -- hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	signal hps_0_h2f_axi_master_bready                                   : std_logic;                      -- hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	signal hps_0_h2f_axi_master_rlast                                    : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	signal hps_0_h2f_axi_master_wlast                                    : std_logic;                      -- hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	signal hps_0_h2f_axi_master_rresp                                    : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	signal hps_0_h2f_axi_master_awid                                     : std_logic_vector(11 downto 0);  -- hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	signal hps_0_h2f_axi_master_bid                                      : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	signal hps_0_h2f_axi_master_bvalid                                   : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	signal hps_0_h2f_axi_master_awsize                                   : std_logic_vector(2 downto 0);   -- hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	signal hps_0_h2f_axi_master_awvalid                                  : std_logic;                      -- hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	signal hps_0_h2f_axi_master_rvalid                                   : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_readdata            : std_logic_vector(63 downto 0);  -- FPGA_Slave_mm_bridge:s0_readdata -> mm_interconnect_1:FPGA_Slave_mm_bridge_s0_readdata
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_waitrequest         : std_logic;                      -- FPGA_Slave_mm_bridge:s0_waitrequest -> mm_interconnect_1:FPGA_Slave_mm_bridge_s0_waitrequest
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_debugaccess         : std_logic;                      -- mm_interconnect_1:FPGA_Slave_mm_bridge_s0_debugaccess -> FPGA_Slave_mm_bridge:s0_debugaccess
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_address             : std_logic_vector(17 downto 0);  -- mm_interconnect_1:FPGA_Slave_mm_bridge_s0_address -> FPGA_Slave_mm_bridge:s0_address
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_read                : std_logic;                      -- mm_interconnect_1:FPGA_Slave_mm_bridge_s0_read -> FPGA_Slave_mm_bridge:s0_read
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_byteenable          : std_logic_vector(7 downto 0);   -- mm_interconnect_1:FPGA_Slave_mm_bridge_s0_byteenable -> FPGA_Slave_mm_bridge:s0_byteenable
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_readdatavalid       : std_logic;                      -- FPGA_Slave_mm_bridge:s0_readdatavalid -> mm_interconnect_1:FPGA_Slave_mm_bridge_s0_readdatavalid
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_write               : std_logic;                      -- mm_interconnect_1:FPGA_Slave_mm_bridge_s0_write -> FPGA_Slave_mm_bridge:s0_write
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_writedata           : std_logic_vector(63 downto 0);  -- mm_interconnect_1:FPGA_Slave_mm_bridge_s0_writedata -> FPGA_Slave_mm_bridge:s0_writedata
	signal mm_interconnect_1_fpga_slave_mm_bridge_s0_burstcount          : std_logic_vector(0 downto 0);   -- mm_interconnect_1:FPGA_Slave_mm_bridge_s0_burstcount -> FPGA_Slave_mm_bridge:s0_burstcount
	signal hps_0_h2f_lw_axi_master_awburst                               : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                                 : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                                 : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_WSTRB -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                                : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                   : std_logic_vector(11 downto 0);  -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                                : std_logic;                      -- hps_0:h2f_lw_RREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                                 : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                   : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_WID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                               : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                                : std_logic;                      -- hps_0:h2f_lw_WVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                                : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_ARADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                                : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                                : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                                 : std_logic_vector(31 downto 0);  -- hps_0:h2f_lw_WDATA -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                               : std_logic;                      -- hps_0:h2f_lw_ARVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                               : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                                  : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_ARID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                                : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                                : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                                : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_AWADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_2:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                               : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                                 : std_logic_vector(31 downto 0);  -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                               : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                               : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                                : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                                : std_logic;                      -- hps_0:h2f_lw_BREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                                 : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                                 : std_logic;                      -- hps_0:h2f_lw_WLAST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                                  : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_AWID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                   : std_logic_vector(11 downto 0);  -- mm_interconnect_2:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                                : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                                : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                               : std_logic;                      -- hps_0:h2f_lw_AWVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                                : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal fpga_only_master_master_readdata                              : std_logic_vector(31 downto 0);  -- mm_interconnect_2:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	signal fpga_only_master_master_waitrequest                           : std_logic;                      -- mm_interconnect_2:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	signal fpga_only_master_master_address                               : std_logic_vector(31 downto 0);  -- fpga_only_master:master_address -> mm_interconnect_2:fpga_only_master_master_address
	signal fpga_only_master_master_read                                  : std_logic;                      -- fpga_only_master:master_read -> mm_interconnect_2:fpga_only_master_master_read
	signal fpga_only_master_master_byteenable                            : std_logic_vector(3 downto 0);   -- fpga_only_master:master_byteenable -> mm_interconnect_2:fpga_only_master_master_byteenable
	signal fpga_only_master_master_readdatavalid                         : std_logic;                      -- mm_interconnect_2:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	signal fpga_only_master_master_write                                 : std_logic;                      -- fpga_only_master:master_write -> mm_interconnect_2:fpga_only_master_master_write
	signal fpga_only_master_master_writedata                             : std_logic_vector(31 downto 0);  -- fpga_only_master:master_writedata -> mm_interconnect_2:fpga_only_master_master_writedata
	signal mm_interconnect_2_lw_mm_bridge_s0_readdata                    : std_logic_vector(31 downto 0);  -- lw_mm_bridge:s0_readdata -> mm_interconnect_2:lw_mm_bridge_s0_readdata
	signal mm_interconnect_2_lw_mm_bridge_s0_waitrequest                 : std_logic;                      -- lw_mm_bridge:s0_waitrequest -> mm_interconnect_2:lw_mm_bridge_s0_waitrequest
	signal mm_interconnect_2_lw_mm_bridge_s0_debugaccess                 : std_logic;                      -- mm_interconnect_2:lw_mm_bridge_s0_debugaccess -> lw_mm_bridge:s0_debugaccess
	signal mm_interconnect_2_lw_mm_bridge_s0_address                     : std_logic_vector(19 downto 0);  -- mm_interconnect_2:lw_mm_bridge_s0_address -> lw_mm_bridge:s0_address
	signal mm_interconnect_2_lw_mm_bridge_s0_read                        : std_logic;                      -- mm_interconnect_2:lw_mm_bridge_s0_read -> lw_mm_bridge:s0_read
	signal mm_interconnect_2_lw_mm_bridge_s0_byteenable                  : std_logic_vector(3 downto 0);   -- mm_interconnect_2:lw_mm_bridge_s0_byteenable -> lw_mm_bridge:s0_byteenable
	signal mm_interconnect_2_lw_mm_bridge_s0_readdatavalid               : std_logic;                      -- lw_mm_bridge:s0_readdatavalid -> mm_interconnect_2:lw_mm_bridge_s0_readdatavalid
	signal mm_interconnect_2_lw_mm_bridge_s0_write                       : std_logic;                      -- mm_interconnect_2:lw_mm_bridge_s0_write -> lw_mm_bridge:s0_write
	signal mm_interconnect_2_lw_mm_bridge_s0_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_2:lw_mm_bridge_s0_writedata -> lw_mm_bridge:s0_writedata
	signal mm_interconnect_2_lw_mm_bridge_s0_burstcount                  : std_logic_vector(0 downto 0);   -- mm_interconnect_2:lw_mm_bridge_s0_burstcount -> lw_mm_bridge:s0_burstcount
	signal lw_mm_bridge_m0_waitrequest                                   : std_logic;                      -- mm_interconnect_3:lw_mm_bridge_m0_waitrequest -> lw_mm_bridge:m0_waitrequest
	signal lw_mm_bridge_m0_readdata                                      : std_logic_vector(31 downto 0);  -- mm_interconnect_3:lw_mm_bridge_m0_readdata -> lw_mm_bridge:m0_readdata
	signal lw_mm_bridge_m0_debugaccess                                   : std_logic;                      -- lw_mm_bridge:m0_debugaccess -> mm_interconnect_3:lw_mm_bridge_m0_debugaccess
	signal lw_mm_bridge_m0_address                                       : std_logic_vector(19 downto 0);  -- lw_mm_bridge:m0_address -> mm_interconnect_3:lw_mm_bridge_m0_address
	signal lw_mm_bridge_m0_read                                          : std_logic;                      -- lw_mm_bridge:m0_read -> mm_interconnect_3:lw_mm_bridge_m0_read
	signal lw_mm_bridge_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- lw_mm_bridge:m0_byteenable -> mm_interconnect_3:lw_mm_bridge_m0_byteenable
	signal lw_mm_bridge_m0_readdatavalid                                 : std_logic;                      -- mm_interconnect_3:lw_mm_bridge_m0_readdatavalid -> lw_mm_bridge:m0_readdatavalid
	signal lw_mm_bridge_m0_writedata                                     : std_logic_vector(31 downto 0);  -- lw_mm_bridge:m0_writedata -> mm_interconnect_3:lw_mm_bridge_m0_writedata
	signal lw_mm_bridge_m0_write                                         : std_logic;                      -- lw_mm_bridge:m0_write -> mm_interconnect_3:lw_mm_bridge_m0_write
	signal lw_mm_bridge_m0_burstcount                                    : std_logic_vector(0 downto 0);   -- lw_mm_bridge:m0_burstcount -> mm_interconnect_3:lw_mm_bridge_m0_burstcount
	signal mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata     : std_logic_vector(31 downto 0);  -- intr_capturer_0:rddata -> mm_interconnect_3:intr_capturer_0_avalon_slave_0_readdata
	signal mm_interconnect_3_intr_capturer_0_avalon_slave_0_address      : std_logic_vector(0 downto 0);   -- mm_interconnect_3:intr_capturer_0_avalon_slave_0_address -> intr_capturer_0:addr
	signal mm_interconnect_3_intr_capturer_0_avalon_slave_0_read         : std_logic;                      -- mm_interconnect_3:intr_capturer_0_avalon_slave_0_read -> intr_capturer_0:read
	signal mm_interconnect_3_sysid_qsys_control_slave_readdata           : std_logic_vector(31 downto 0);  -- sysid_qsys:readdata -> mm_interconnect_3:sysid_qsys_control_slave_readdata
	signal mm_interconnect_3_sysid_qsys_control_slave_address            : std_logic_vector(0 downto 0);   -- mm_interconnect_3:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_3_kbandipsub_slw_readdata                     : std_logic_vector(31 downto 0);  -- KBandIPsub:slw_readdata -> mm_interconnect_3:KBandIPsub_slw_readdata
	signal mm_interconnect_3_kbandipsub_slw_waitrequest                  : std_logic;                      -- KBandIPsub:slw_waitrequest -> mm_interconnect_3:KBandIPsub_slw_waitrequest
	signal mm_interconnect_3_kbandipsub_slw_debugaccess                  : std_logic;                      -- mm_interconnect_3:KBandIPsub_slw_debugaccess -> KBandIPsub:slw_debugaccess
	signal mm_interconnect_3_kbandipsub_slw_address                      : std_logic_vector(16 downto 0);  -- mm_interconnect_3:KBandIPsub_slw_address -> KBandIPsub:slw_address
	signal mm_interconnect_3_kbandipsub_slw_read                         : std_logic;                      -- mm_interconnect_3:KBandIPsub_slw_read -> KBandIPsub:slw_read
	signal mm_interconnect_3_kbandipsub_slw_byteenable                   : std_logic_vector(3 downto 0);   -- mm_interconnect_3:KBandIPsub_slw_byteenable -> KBandIPsub:slw_byteenable
	signal mm_interconnect_3_kbandipsub_slw_readdatavalid                : std_logic;                      -- KBandIPsub:slw_readdatavalid -> mm_interconnect_3:KBandIPsub_slw_readdatavalid
	signal mm_interconnect_3_kbandipsub_slw_write                        : std_logic;                      -- mm_interconnect_3:KBandIPsub_slw_write -> KBandIPsub:slw_write
	signal mm_interconnect_3_kbandipsub_slw_writedata                    : std_logic_vector(31 downto 0);  -- mm_interconnect_3:KBandIPsub_slw_writedata -> KBandIPsub:slw_writedata
	signal mm_interconnect_3_kbandipsub_slw_burstcount                   : std_logic_vector(0 downto 0);   -- mm_interconnect_3:KBandIPsub_slw_burstcount -> KBandIPsub:slw_burstcount
	signal kbandipsub_m0_waitrequest                                     : std_logic;                      -- mm_interconnect_6:KBandIPsub_m0_waitrequest -> KBandIPsub:m0_waitrequest
	signal kbandipsub_m0_readdata                                        : std_logic_vector(127 downto 0); -- mm_interconnect_6:KBandIPsub_m0_readdata -> KBandIPsub:m0_readdata
	signal kbandipsub_m0_debugaccess                                     : std_logic;                      -- KBandIPsub:m0_debugaccess -> mm_interconnect_6:KBandIPsub_m0_debugaccess
	signal kbandipsub_m0_address                                         : std_logic_vector(29 downto 0);  -- KBandIPsub:m0_address -> mm_interconnect_6:KBandIPsub_m0_address
	signal kbandipsub_m0_read                                            : std_logic;                      -- KBandIPsub:m0_read -> mm_interconnect_6:KBandIPsub_m0_read
	signal kbandipsub_m0_byteenable                                      : std_logic_vector(15 downto 0);  -- KBandIPsub:m0_byteenable -> mm_interconnect_6:KBandIPsub_m0_byteenable
	signal kbandipsub_m0_readdatavalid                                   : std_logic;                      -- mm_interconnect_6:KBandIPsub_m0_readdatavalid -> KBandIPsub:m0_readdatavalid
	signal kbandipsub_m0_writedata                                       : std_logic_vector(127 downto 0); -- KBandIPsub:m0_writedata -> mm_interconnect_6:KBandIPsub_m0_writedata
	signal kbandipsub_m0_write                                           : std_logic;                      -- KBandIPsub:m0_write -> mm_interconnect_6:KBandIPsub_m0_write
	signal kbandipsub_m0_burstcount                                      : std_logic_vector(4 downto 0);   -- KBandIPsub:m0_burstcount -> mm_interconnect_6:KBandIPsub_m0_burstcount
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdata      : std_logic_vector(127 downto 0); -- fft_ddr_bridge:avs_s0_readdata -> mm_interconnect_6:fft_ddr_bridge_windowed_slave_readdata
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_waitrequest   : std_logic;                      -- fft_ddr_bridge:avs_s0_waitrequest -> mm_interconnect_6:fft_ddr_bridge_windowed_slave_waitrequest
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_address       : std_logic_vector(25 downto 0);  -- mm_interconnect_6:fft_ddr_bridge_windowed_slave_address -> fft_ddr_bridge:avs_s0_address
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_read          : std_logic;                      -- mm_interconnect_6:fft_ddr_bridge_windowed_slave_read -> fft_ddr_bridge:avs_s0_read
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_byteenable    : std_logic_vector(15 downto 0);  -- mm_interconnect_6:fft_ddr_bridge_windowed_slave_byteenable -> fft_ddr_bridge:avs_s0_byteenable
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdatavalid : std_logic;                      -- fft_ddr_bridge:avs_s0_readdatavalid -> mm_interconnect_6:fft_ddr_bridge_windowed_slave_readdatavalid
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_write         : std_logic;                      -- mm_interconnect_6:fft_ddr_bridge_windowed_slave_write -> fft_ddr_bridge:avs_s0_write
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_writedata     : std_logic_vector(127 downto 0); -- mm_interconnect_6:fft_ddr_bridge_windowed_slave_writedata -> fft_ddr_bridge:avs_s0_writedata
	signal mm_interconnect_6_fft_ddr_bridge_windowed_slave_burstcount    : std_logic_vector(4 downto 0);   -- mm_interconnect_6:fft_ddr_bridge_windowed_slave_burstcount -> fft_ddr_bridge:avs_s0_burstcount
	signal hps_0_f2h_irq0_irq                                            : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	signal hps_0_f2h_irq1_irq                                            : std_logic_vector(31 downto 0);  -- irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	signal intr_capturer_0_interrupt_receiver_irq                        : std_logic_vector(31 downto 0);  -- irq_mapper_002:sender_irq -> intr_capturer_0:interrupt_in
	signal irq_mapper_receiver0_irq                                      : std_logic;                      -- KBandIPsub:kbandinput_1_csr_irq_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver0_irq]
	signal irq_mapper_receiver1_irq                                      : std_logic;                      -- KBandIPsub:kbandinput_2_csr_irq_irq -> [irq_mapper:receiver1_irq, irq_mapper_002:receiver1_irq]
	signal irq_mapper_receiver2_irq                                      : std_logic;                      -- KBandIPsub:kbandoutput_csr_irq_irq -> [irq_mapper:receiver2_irq, irq_mapper_002:receiver2_irq]
	signal rst_controller_reset_out_reset                                : std_logic;                      -- rst_controller:reset_out -> [FPGA_Slave_mm_bridge:reset, axi_bridge_for_acp_128_0:reset, fft_ddr_bridge:reset, irq_mapper_002:reset, lw_mm_bridge:reset, mm_interconnect_0:fft_ddr_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:FPGA_Slave_mm_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_2:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:lw_mm_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_3:KBandIPsub_reset_reset_bridge_in_reset_reset, mm_interconnect_3:lw_mm_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_6:KBandIPsub_reset_reset_bridge_in_reset_reset, mm_interconnect_6:fft_ddr_bridge_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                      -- rst_controller_001:reset_out -> [mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                       : std_logic;                      -- reset_reset_n:inv -> [fpga_only_master:clk_reset_reset, pll_0:rst, rst_controller:reset_in0]
	signal hps_0_h2f_reset_reset_n_ports_inv                             : std_logic;                      -- hps_0_h2f_reset_reset_n:inv -> rst_controller_001:reset_in0
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                      -- rst_controller_reset_out_reset:inv -> [intr_capturer_0:rst_n, sysid_qsys:reset_n]

begin

	fpga_slave_mm_bridge : component soc_system_fpga_slave_mm_bridge
		generic map (
			DATA_WIDTH        => 64,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 18,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => pll_0_outclk0_clk,                                       --   clk.clk
			reset            => rst_controller_reset_out_reset,                          -- reset.reset
			s0_waitrequest   => mm_interconnect_1_fpga_slave_mm_bridge_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_interconnect_1_fpga_slave_mm_bridge_s0_readdata,      --      .readdata
			s0_readdatavalid => mm_interconnect_1_fpga_slave_mm_bridge_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_interconnect_1_fpga_slave_mm_bridge_s0_burstcount,    --      .burstcount
			s0_writedata     => mm_interconnect_1_fpga_slave_mm_bridge_s0_writedata,     --      .writedata
			s0_address       => mm_interconnect_1_fpga_slave_mm_bridge_s0_address,       --      .address
			s0_write         => mm_interconnect_1_fpga_slave_mm_bridge_s0_write,         --      .write
			s0_read          => mm_interconnect_1_fpga_slave_mm_bridge_s0_read,          --      .read
			s0_byteenable    => mm_interconnect_1_fpga_slave_mm_bridge_s0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_interconnect_1_fpga_slave_mm_bridge_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => fpga_slave_mm_bridge_m0_waitrequest,                     --    m0.waitrequest
			m0_readdata      => fpga_slave_mm_bridge_m0_readdata,                        --      .readdata
			m0_readdatavalid => fpga_slave_mm_bridge_m0_readdatavalid,                   --      .readdatavalid
			m0_burstcount    => fpga_slave_mm_bridge_m0_burstcount,                      --      .burstcount
			m0_writedata     => fpga_slave_mm_bridge_m0_writedata,                       --      .writedata
			m0_address       => fpga_slave_mm_bridge_m0_address,                         --      .address
			m0_write         => fpga_slave_mm_bridge_m0_write,                           --      .write
			m0_read          => fpga_slave_mm_bridge_m0_read,                            --      .read
			m0_byteenable    => fpga_slave_mm_bridge_m0_byteenable,                      --      .byteenable
			m0_debugaccess   => fpga_slave_mm_bridge_m0_debugaccess,                     --      .debugaccess
			s0_response      => open,                                                    -- (terminated)
			m0_response      => "00"                                                     -- (terminated)
		);

	kbandipsub : component soc_system_KBandIPsub
		port map (
			clk_clk                  => pll_0_outclk0_clk,                              --                  clk.clk
			clk_int_clk              => pll_0_outclk1_clk,                              --              clk_int.clk
			kbandinput_1_csr_irq_irq => irq_mapper_receiver0_irq,                       -- kbandinput_1_csr_irq.irq
			kbandinput_2_csr_irq_irq => irq_mapper_receiver1_irq,                       -- kbandinput_2_csr_irq.irq
			kbandoutput_csr_irq_irq  => irq_mapper_receiver2_irq,                       --  kbandoutput_csr_irq.irq
			m0_waitrequest           => kbandipsub_m0_waitrequest,                      --                   m0.waitrequest
			m0_readdata              => kbandipsub_m0_readdata,                         --                     .readdata
			m0_readdatavalid         => kbandipsub_m0_readdatavalid,                    --                     .readdatavalid
			m0_burstcount            => kbandipsub_m0_burstcount,                       --                     .burstcount
			m0_writedata             => kbandipsub_m0_writedata,                        --                     .writedata
			m0_address               => kbandipsub_m0_address,                          --                     .address
			m0_write                 => kbandipsub_m0_write,                            --                     .write
			m0_read                  => kbandipsub_m0_read,                             --                     .read
			m0_byteenable            => kbandipsub_m0_byteenable,                       --                     .byteenable
			m0_debugaccess           => kbandipsub_m0_debugaccess,                      --                     .debugaccess
			reset_reset_n            => reset_reset_n,                                  --                reset.reset_n
			sfpga_waitrequest        => fpga_slave_mm_bridge_m0_waitrequest,            --                sfpga.waitrequest
			sfpga_readdata           => fpga_slave_mm_bridge_m0_readdata,               --                     .readdata
			sfpga_readdatavalid      => fpga_slave_mm_bridge_m0_readdatavalid,          --                     .readdatavalid
			sfpga_burstcount         => fpga_slave_mm_bridge_m0_burstcount,             --                     .burstcount
			sfpga_writedata          => fpga_slave_mm_bridge_m0_writedata,              --                     .writedata
			sfpga_address            => fpga_slave_mm_bridge_m0_address,                --                     .address
			sfpga_write              => fpga_slave_mm_bridge_m0_write,                  --                     .write
			sfpga_read               => fpga_slave_mm_bridge_m0_read,                   --                     .read
			sfpga_byteenable         => fpga_slave_mm_bridge_m0_byteenable,             --                     .byteenable
			sfpga_debugaccess        => fpga_slave_mm_bridge_m0_debugaccess,            --                     .debugaccess
			slw_waitrequest          => mm_interconnect_3_kbandipsub_slw_waitrequest,   --                  slw.waitrequest
			slw_readdata             => mm_interconnect_3_kbandipsub_slw_readdata,      --                     .readdata
			slw_readdatavalid        => mm_interconnect_3_kbandipsub_slw_readdatavalid, --                     .readdatavalid
			slw_burstcount           => mm_interconnect_3_kbandipsub_slw_burstcount,    --                     .burstcount
			slw_writedata            => mm_interconnect_3_kbandipsub_slw_writedata,     --                     .writedata
			slw_address              => mm_interconnect_3_kbandipsub_slw_address,       --                     .address
			slw_write                => mm_interconnect_3_kbandipsub_slw_write,         --                     .write
			slw_read                 => mm_interconnect_3_kbandipsub_slw_read,          --                     .read
			slw_byteenable           => mm_interconnect_3_kbandipsub_slw_byteenable,    --                     .byteenable
			slw_debugaccess          => mm_interconnect_3_kbandipsub_slw_debugaccess    --                     .debugaccess
		);

	axi_bridge_for_acp_128_0 : component axi_bridge_for_acp_128
		port map (
			clk            => pll_0_outclk0_clk,                                     -- clock.clk
			reset          => rst_controller_reset_out_reset,                        -- reset.reset
			axm_m0_araddr  => axi_bridge_for_acp_128_0_m0_araddr,                    --    m0.araddr
			axm_m0_arburst => axi_bridge_for_acp_128_0_m0_arburst,                   --      .arburst
			axm_m0_arcache => axi_bridge_for_acp_128_0_m0_arcache,                   --      .arcache
			axm_m0_arid    => axi_bridge_for_acp_128_0_m0_arid,                      --      .arid
			axm_m0_arlen   => axi_bridge_for_acp_128_0_m0_arlen,                     --      .arlen
			axm_m0_arlock  => axi_bridge_for_acp_128_0_m0_arlock,                    --      .arlock
			axm_m0_arprot  => axi_bridge_for_acp_128_0_m0_arprot,                    --      .arprot
			axm_m0_arready => axi_bridge_for_acp_128_0_m0_arready,                   --      .arready
			axm_m0_arsize  => axi_bridge_for_acp_128_0_m0_arsize,                    --      .arsize
			axm_m0_aruser  => axi_bridge_for_acp_128_0_m0_aruser,                    --      .aruser
			axm_m0_arvalid => axi_bridge_for_acp_128_0_m0_arvalid,                   --      .arvalid
			axm_m0_awaddr  => axi_bridge_for_acp_128_0_m0_awaddr,                    --      .awaddr
			axm_m0_awburst => axi_bridge_for_acp_128_0_m0_awburst,                   --      .awburst
			axm_m0_awcache => axi_bridge_for_acp_128_0_m0_awcache,                   --      .awcache
			axm_m0_awid    => axi_bridge_for_acp_128_0_m0_awid,                      --      .awid
			axm_m0_awlen   => axi_bridge_for_acp_128_0_m0_awlen,                     --      .awlen
			axm_m0_awlock  => axi_bridge_for_acp_128_0_m0_awlock,                    --      .awlock
			axm_m0_awprot  => axi_bridge_for_acp_128_0_m0_awprot,                    --      .awprot
			axm_m0_awready => axi_bridge_for_acp_128_0_m0_awready,                   --      .awready
			axm_m0_awsize  => axi_bridge_for_acp_128_0_m0_awsize,                    --      .awsize
			axm_m0_awuser  => axi_bridge_for_acp_128_0_m0_awuser,                    --      .awuser
			axm_m0_awvalid => axi_bridge_for_acp_128_0_m0_awvalid,                   --      .awvalid
			axm_m0_bid     => axi_bridge_for_acp_128_0_m0_bid,                       --      .bid
			axm_m0_bready  => axi_bridge_for_acp_128_0_m0_bready,                    --      .bready
			axm_m0_bresp   => axi_bridge_for_acp_128_0_m0_bresp,                     --      .bresp
			axm_m0_bvalid  => axi_bridge_for_acp_128_0_m0_bvalid,                    --      .bvalid
			axm_m0_rdata   => axi_bridge_for_acp_128_0_m0_rdata,                     --      .rdata
			axm_m0_rid     => axi_bridge_for_acp_128_0_m0_rid,                       --      .rid
			axm_m0_rlast   => axi_bridge_for_acp_128_0_m0_rlast,                     --      .rlast
			axm_m0_rready  => axi_bridge_for_acp_128_0_m0_rready,                    --      .rready
			axm_m0_rresp   => axi_bridge_for_acp_128_0_m0_rresp,                     --      .rresp
			axm_m0_rvalid  => axi_bridge_for_acp_128_0_m0_rvalid,                    --      .rvalid
			axm_m0_wdata   => axi_bridge_for_acp_128_0_m0_wdata,                     --      .wdata
			axm_m0_wid     => axi_bridge_for_acp_128_0_m0_wid,                       --      .wid
			axm_m0_wlast   => axi_bridge_for_acp_128_0_m0_wlast,                     --      .wlast
			axm_m0_wready  => axi_bridge_for_acp_128_0_m0_wready,                    --      .wready
			axm_m0_wstrb   => axi_bridge_for_acp_128_0_m0_wstrb,                     --      .wstrb
			axm_m0_wvalid  => axi_bridge_for_acp_128_0_m0_wvalid,                    --      .wvalid
			axs_s0_araddr  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_araddr,  --    s0.araddr
			axs_s0_arburst => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arburst, --      .arburst
			axs_s0_arcache => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arcache, --      .arcache
			axs_s0_arid    => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arid,    --      .arid
			axs_s0_arlen   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlen,   --      .arlen
			axs_s0_arlock  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlock,  --      .arlock
			axs_s0_arprot  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arprot,  --      .arprot
			axs_s0_arready => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arready, --      .arready
			axs_s0_arsize  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arsize,  --      .arsize
			axs_s0_aruser  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_aruser,  --      .aruser
			axs_s0_arvalid => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arvalid, --      .arvalid
			axs_s0_awaddr  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awaddr,  --      .awaddr
			axs_s0_awburst => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awburst, --      .awburst
			axs_s0_awcache => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awcache, --      .awcache
			axs_s0_awid    => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awid,    --      .awid
			axs_s0_awlen   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlen,   --      .awlen
			axs_s0_awlock  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlock,  --      .awlock
			axs_s0_awprot  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awprot,  --      .awprot
			axs_s0_awready => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awready, --      .awready
			axs_s0_awsize  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awsize,  --      .awsize
			axs_s0_awuser  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awuser,  --      .awuser
			axs_s0_awvalid => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awvalid, --      .awvalid
			axs_s0_bid     => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bid,     --      .bid
			axs_s0_bready  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bready,  --      .bready
			axs_s0_bresp   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bresp,   --      .bresp
			axs_s0_bvalid  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bvalid,  --      .bvalid
			axs_s0_rdata   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rdata,   --      .rdata
			axs_s0_rid     => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rid,     --      .rid
			axs_s0_rlast   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rlast,   --      .rlast
			axs_s0_rready  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rready,  --      .rready
			axs_s0_rresp   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rresp,   --      .rresp
			axs_s0_rvalid  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rvalid,  --      .rvalid
			axs_s0_wdata   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wdata,   --      .wdata
			axs_s0_wid     => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wid,     --      .wid
			axs_s0_wlast   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wlast,   --      .wlast
			axs_s0_wready  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wready,  --      .wready
			axs_s0_wstrb   => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wstrb,   --      .wstrb
			axs_s0_wvalid  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wvalid   --      .wvalid
		);

	fft_ddr_bridge : component altera_address_span_extender
		generic map (
			DATA_WIDTH           => 128,
			BYTEENABLE_WIDTH     => 16,
			MASTER_ADDRESS_WIDTH => 32,
			SLAVE_ADDRESS_WIDTH  => 26,
			SLAVE_ADDRESS_SHIFT  => 4,
			BURSTCOUNT_WIDTH     => 5,
			CNTL_ADDRESS_WIDTH   => 1,
			SUB_WINDOW_COUNT     => 1,
			MASTER_ADDRESS_DEF   => "0000000000000000000000000000000010000000000000000000000000000000"
		)
		port map (
			clk                  => pll_0_outclk0_clk,                                             --           clock.clk
			reset                => rst_controller_reset_out_reset,                                --           reset.reset
			avs_s0_address       => mm_interconnect_6_fft_ddr_bridge_windowed_slave_address,       --  windowed_slave.address
			avs_s0_read          => mm_interconnect_6_fft_ddr_bridge_windowed_slave_read,          --                .read
			avs_s0_readdata      => mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdata,      --                .readdata
			avs_s0_write         => mm_interconnect_6_fft_ddr_bridge_windowed_slave_write,         --                .write
			avs_s0_writedata     => mm_interconnect_6_fft_ddr_bridge_windowed_slave_writedata,     --                .writedata
			avs_s0_readdatavalid => mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdatavalid, --                .readdatavalid
			avs_s0_waitrequest   => mm_interconnect_6_fft_ddr_bridge_windowed_slave_waitrequest,   --                .waitrequest
			avs_s0_byteenable    => mm_interconnect_6_fft_ddr_bridge_windowed_slave_byteenable,    --                .byteenable
			avs_s0_burstcount    => mm_interconnect_6_fft_ddr_bridge_windowed_slave_burstcount,    --                .burstcount
			avm_m0_address       => fft_ddr_bridge_expanded_master_address,                        -- expanded_master.address
			avm_m0_read          => fft_ddr_bridge_expanded_master_read,                           --                .read
			avm_m0_waitrequest   => fft_ddr_bridge_expanded_master_waitrequest,                    --                .waitrequest
			avm_m0_readdata      => fft_ddr_bridge_expanded_master_readdata,                       --                .readdata
			avm_m0_write         => fft_ddr_bridge_expanded_master_write,                          --                .write
			avm_m0_writedata     => fft_ddr_bridge_expanded_master_writedata,                      --                .writedata
			avm_m0_readdatavalid => fft_ddr_bridge_expanded_master_readdatavalid,                  --                .readdatavalid
			avm_m0_byteenable    => fft_ddr_bridge_expanded_master_byteenable,                     --                .byteenable
			avm_m0_burstcount    => fft_ddr_bridge_expanded_master_burstcount,                     --                .burstcount
			avs_cntl_read        => open,                                                          --            cntl.read
			avs_cntl_readdata    => open,                                                          --                .readdata
			avs_cntl_write       => open,                                                          --                .write
			avs_cntl_writedata   => open,                                                          --                .writedata
			avs_cntl_byteenable  => open,                                                          --                .byteenable
			avs_cntl_address     => "0"                                                            --     (terminated)
		);

	fpga_only_master : component soc_system_fpga_only_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => pll_0_outclk0_clk,                     --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,               --    clk_reset.reset
			master_address       => fpga_only_master_master_address,       --       master.address
			master_readdata      => fpga_only_master_master_readdata,      --             .readdata
			master_read          => fpga_only_master_master_read,          --             .read
			master_write         => fpga_only_master_master_write,         --             .write
			master_writedata     => fpga_only_master_master_writedata,     --             .writedata
			master_waitrequest   => fpga_only_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => fpga_only_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => fpga_only_master_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                   -- master_reset.reset
		);

	hps_0 : component soc_system_hps_0
		generic map (
			F2S_Width => 3,
			S2F_Width => 2
		)
		port map (
			f2h_cold_rst_req_n       => hps_0_f2h_cold_reset_req_reset_n,      --  f2h_cold_reset_req.reset_n
			f2h_dbg_rst_req_n        => hps_0_f2h_debug_reset_req_reset_n,     -- f2h_debug_reset_req.reset_n
			f2h_warm_rst_req_n       => hps_0_f2h_warm_reset_req_reset_n,      --  f2h_warm_reset_req.reset_n
			h2f_user0_clk            => open,                                  --     h2f_user0_clock.clk
			h2f_user1_clk            => open,                                  --     h2f_user1_clock.clk
			f2h_stm_hwevents         => hps_0_f2h_stm_hw_events_stm_hwevents,  --   f2h_stm_hw_events.stm_hwevents
			mem_a                    => memory_mem_a,                          --              memory.mem_a
			mem_ba                   => memory_mem_ba,                         --                    .mem_ba
			mem_ck                   => memory_mem_ck,                         --                    .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                       --                    .mem_ck_n
			mem_cke                  => memory_mem_cke,                        --                    .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                       --                    .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                      --                    .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                      --                    .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                       --                    .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                    --                    .mem_reset_n
			mem_dq                   => memory_mem_dq,                         --                    .mem_dq
			mem_dqs                  => memory_mem_dqs,                        --                    .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                      --                    .mem_dqs_n
			mem_odt                  => memory_mem_odt,                        --                    .mem_odt
			mem_dm                   => memory_mem_dm,                         --                    .mem_dm
			oct_rzqin                => memory_oct_rzqin,                      --                    .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_0_hps_io_hps_io_emac1_inst_TX_CLK, --              hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_0_hps_io_hps_io_emac1_inst_TXD0,   --                    .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_0_hps_io_hps_io_emac1_inst_TXD1,   --                    .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_0_hps_io_hps_io_emac1_inst_TXD2,   --                    .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_0_hps_io_hps_io_emac1_inst_TXD3,   --                    .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_0_hps_io_hps_io_emac1_inst_RXD0,   --                    .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_0_hps_io_hps_io_emac1_inst_MDIO,   --                    .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_0_hps_io_hps_io_emac1_inst_MDC,    --                    .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_0_hps_io_hps_io_emac1_inst_RX_CTL, --                    .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_0_hps_io_hps_io_emac1_inst_TX_CTL, --                    .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_0_hps_io_hps_io_emac1_inst_RX_CLK, --                    .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_0_hps_io_hps_io_emac1_inst_RXD1,   --                    .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_0_hps_io_hps_io_emac1_inst_RXD2,   --                    .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_0_hps_io_hps_io_emac1_inst_RXD3,   --                    .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_0_hps_io_hps_io_sdio_inst_CMD,     --                    .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_0_hps_io_hps_io_sdio_inst_D0,      --                    .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_0_hps_io_hps_io_sdio_inst_D1,      --                    .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_0_hps_io_hps_io_sdio_inst_CLK,     --                    .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_0_hps_io_hps_io_sdio_inst_D2,      --                    .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_0_hps_io_hps_io_sdio_inst_D3,      --                    .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_0_hps_io_hps_io_usb1_inst_D0,      --                    .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_0_hps_io_hps_io_usb1_inst_D1,      --                    .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_0_hps_io_hps_io_usb1_inst_D2,      --                    .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_0_hps_io_hps_io_usb1_inst_D3,      --                    .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_0_hps_io_hps_io_usb1_inst_D4,      --                    .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_0_hps_io_hps_io_usb1_inst_D5,      --                    .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_0_hps_io_hps_io_usb1_inst_D6,      --                    .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_0_hps_io_hps_io_usb1_inst_D7,      --                    .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_0_hps_io_hps_io_usb1_inst_CLK,     --                    .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_0_hps_io_hps_io_usb1_inst_STP,     --                    .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_0_hps_io_hps_io_usb1_inst_DIR,     --                    .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_0_hps_io_hps_io_usb1_inst_NXT,     --                    .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_0_hps_io_hps_io_spim1_inst_CLK,    --                    .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_0_hps_io_hps_io_spim1_inst_MOSI,   --                    .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_0_hps_io_hps_io_spim1_inst_MISO,   --                    .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_0_hps_io_hps_io_spim1_inst_SS0,    --                    .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_0_hps_io_hps_io_uart0_inst_RX,     --                    .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_0_hps_io_hps_io_uart0_inst_TX,     --                    .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_0_hps_io_hps_io_i2c0_inst_SDA,     --                    .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_0_hps_io_hps_io_i2c0_inst_SCL,     --                    .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_0_hps_io_hps_io_i2c1_inst_SDA,     --                    .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_0_hps_io_hps_io_i2c1_inst_SCL,     --                    .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_0_hps_io_hps_io_gpio_inst_GPIO09,  --                    .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_0_hps_io_hps_io_gpio_inst_GPIO35,  --                    .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_0_hps_io_hps_io_gpio_inst_GPIO40,  --                    .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  => hps_0_hps_io_hps_io_gpio_inst_GPIO53,  --                    .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_0_hps_io_hps_io_gpio_inst_GPIO54,  --                    .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_0_hps_io_hps_io_gpio_inst_GPIO61,  --                    .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_0_h2f_reset_reset,                 --           h2f_reset.reset_n
			f2h_sdram0_clk           => pll_0_outclk0_clk,                     --    f2h_sdram0_clock.clk
			f2h_sdram0_ADDRESS       => open,                                  --     f2h_sdram0_data.address
			f2h_sdram0_BURSTCOUNT    => open,                                  --                    .burstcount
			f2h_sdram0_WAITREQUEST   => open,                                  --                    .waitrequest
			f2h_sdram0_READDATA      => open,                                  --                    .readdata
			f2h_sdram0_READDATAVALID => open,                                  --                    .readdatavalid
			f2h_sdram0_READ          => open,                                  --                    .read
			f2h_sdram0_WRITEDATA     => open,                                  --                    .writedata
			f2h_sdram0_BYTEENABLE    => open,                                  --                    .byteenable
			f2h_sdram0_WRITE         => open,                                  --                    .write
			h2f_axi_clk              => pll_0_outclk0_clk,                     --       h2f_axi_clock.clk
			h2f_AWID                 => hps_0_h2f_axi_master_awid,             --      h2f_axi_master.awid
			h2f_AWADDR               => hps_0_h2f_axi_master_awaddr,           --                    .awaddr
			h2f_AWLEN                => hps_0_h2f_axi_master_awlen,            --                    .awlen
			h2f_AWSIZE               => hps_0_h2f_axi_master_awsize,           --                    .awsize
			h2f_AWBURST              => hps_0_h2f_axi_master_awburst,          --                    .awburst
			h2f_AWLOCK               => hps_0_h2f_axi_master_awlock,           --                    .awlock
			h2f_AWCACHE              => hps_0_h2f_axi_master_awcache,          --                    .awcache
			h2f_AWPROT               => hps_0_h2f_axi_master_awprot,           --                    .awprot
			h2f_AWVALID              => hps_0_h2f_axi_master_awvalid,          --                    .awvalid
			h2f_AWREADY              => hps_0_h2f_axi_master_awready,          --                    .awready
			h2f_WID                  => hps_0_h2f_axi_master_wid,              --                    .wid
			h2f_WDATA                => hps_0_h2f_axi_master_wdata,            --                    .wdata
			h2f_WSTRB                => hps_0_h2f_axi_master_wstrb,            --                    .wstrb
			h2f_WLAST                => hps_0_h2f_axi_master_wlast,            --                    .wlast
			h2f_WVALID               => hps_0_h2f_axi_master_wvalid,           --                    .wvalid
			h2f_WREADY               => hps_0_h2f_axi_master_wready,           --                    .wready
			h2f_BID                  => hps_0_h2f_axi_master_bid,              --                    .bid
			h2f_BRESP                => hps_0_h2f_axi_master_bresp,            --                    .bresp
			h2f_BVALID               => hps_0_h2f_axi_master_bvalid,           --                    .bvalid
			h2f_BREADY               => hps_0_h2f_axi_master_bready,           --                    .bready
			h2f_ARID                 => hps_0_h2f_axi_master_arid,             --                    .arid
			h2f_ARADDR               => hps_0_h2f_axi_master_araddr,           --                    .araddr
			h2f_ARLEN                => hps_0_h2f_axi_master_arlen,            --                    .arlen
			h2f_ARSIZE               => hps_0_h2f_axi_master_arsize,           --                    .arsize
			h2f_ARBURST              => hps_0_h2f_axi_master_arburst,          --                    .arburst
			h2f_ARLOCK               => hps_0_h2f_axi_master_arlock,           --                    .arlock
			h2f_ARCACHE              => hps_0_h2f_axi_master_arcache,          --                    .arcache
			h2f_ARPROT               => hps_0_h2f_axi_master_arprot,           --                    .arprot
			h2f_ARVALID              => hps_0_h2f_axi_master_arvalid,          --                    .arvalid
			h2f_ARREADY              => hps_0_h2f_axi_master_arready,          --                    .arready
			h2f_RID                  => hps_0_h2f_axi_master_rid,              --                    .rid
			h2f_RDATA                => hps_0_h2f_axi_master_rdata,            --                    .rdata
			h2f_RRESP                => hps_0_h2f_axi_master_rresp,            --                    .rresp
			h2f_RLAST                => hps_0_h2f_axi_master_rlast,            --                    .rlast
			h2f_RVALID               => hps_0_h2f_axi_master_rvalid,           --                    .rvalid
			h2f_RREADY               => hps_0_h2f_axi_master_rready,           --                    .rready
			f2h_axi_clk              => pll_0_outclk0_clk,                     --       f2h_axi_clock.clk
			f2h_AWID                 => axi_bridge_for_acp_128_0_m0_awid,      --       f2h_axi_slave.awid
			f2h_AWADDR               => axi_bridge_for_acp_128_0_m0_awaddr,    --                    .awaddr
			f2h_AWLEN                => axi_bridge_for_acp_128_0_m0_awlen,     --                    .awlen
			f2h_AWSIZE               => axi_bridge_for_acp_128_0_m0_awsize,    --                    .awsize
			f2h_AWBURST              => axi_bridge_for_acp_128_0_m0_awburst,   --                    .awburst
			f2h_AWLOCK               => axi_bridge_for_acp_128_0_m0_awlock,    --                    .awlock
			f2h_AWCACHE              => axi_bridge_for_acp_128_0_m0_awcache,   --                    .awcache
			f2h_AWPROT               => axi_bridge_for_acp_128_0_m0_awprot,    --                    .awprot
			f2h_AWVALID              => axi_bridge_for_acp_128_0_m0_awvalid,   --                    .awvalid
			f2h_AWREADY              => axi_bridge_for_acp_128_0_m0_awready,   --                    .awready
			f2h_AWUSER               => axi_bridge_for_acp_128_0_m0_awuser,    --                    .awuser
			f2h_WID                  => axi_bridge_for_acp_128_0_m0_wid,       --                    .wid
			f2h_WDATA                => axi_bridge_for_acp_128_0_m0_wdata,     --                    .wdata
			f2h_WSTRB                => axi_bridge_for_acp_128_0_m0_wstrb,     --                    .wstrb
			f2h_WLAST                => axi_bridge_for_acp_128_0_m0_wlast,     --                    .wlast
			f2h_WVALID               => axi_bridge_for_acp_128_0_m0_wvalid,    --                    .wvalid
			f2h_WREADY               => axi_bridge_for_acp_128_0_m0_wready,    --                    .wready
			f2h_BID                  => axi_bridge_for_acp_128_0_m0_bid,       --                    .bid
			f2h_BRESP                => axi_bridge_for_acp_128_0_m0_bresp,     --                    .bresp
			f2h_BVALID               => axi_bridge_for_acp_128_0_m0_bvalid,    --                    .bvalid
			f2h_BREADY               => axi_bridge_for_acp_128_0_m0_bready,    --                    .bready
			f2h_ARID                 => axi_bridge_for_acp_128_0_m0_arid,      --                    .arid
			f2h_ARADDR               => axi_bridge_for_acp_128_0_m0_araddr,    --                    .araddr
			f2h_ARLEN                => axi_bridge_for_acp_128_0_m0_arlen,     --                    .arlen
			f2h_ARSIZE               => axi_bridge_for_acp_128_0_m0_arsize,    --                    .arsize
			f2h_ARBURST              => axi_bridge_for_acp_128_0_m0_arburst,   --                    .arburst
			f2h_ARLOCK               => axi_bridge_for_acp_128_0_m0_arlock,    --                    .arlock
			f2h_ARCACHE              => axi_bridge_for_acp_128_0_m0_arcache,   --                    .arcache
			f2h_ARPROT               => axi_bridge_for_acp_128_0_m0_arprot,    --                    .arprot
			f2h_ARVALID              => axi_bridge_for_acp_128_0_m0_arvalid,   --                    .arvalid
			f2h_ARREADY              => axi_bridge_for_acp_128_0_m0_arready,   --                    .arready
			f2h_ARUSER               => axi_bridge_for_acp_128_0_m0_aruser,    --                    .aruser
			f2h_RID                  => axi_bridge_for_acp_128_0_m0_rid,       --                    .rid
			f2h_RDATA                => axi_bridge_for_acp_128_0_m0_rdata,     --                    .rdata
			f2h_RRESP                => axi_bridge_for_acp_128_0_m0_rresp,     --                    .rresp
			f2h_RLAST                => axi_bridge_for_acp_128_0_m0_rlast,     --                    .rlast
			f2h_RVALID               => axi_bridge_for_acp_128_0_m0_rvalid,    --                    .rvalid
			f2h_RREADY               => axi_bridge_for_acp_128_0_m0_rready,    --                    .rready
			h2f_lw_axi_clk           => pll_0_outclk0_clk,                     --    h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,          --   h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,        --                    .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,         --                    .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,        --                    .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst,       --                    .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,        --                    .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache,       --                    .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,        --                    .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid,       --                    .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready,       --                    .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,           --                    .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,         --                    .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,         --                    .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,         --                    .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,        --                    .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,        --                    .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,           --                    .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,         --                    .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,        --                    .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,        --                    .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,          --                    .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,        --                    .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,         --                    .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,        --                    .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst,       --                    .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,        --                    .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache,       --                    .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,        --                    .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid,       --                    .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready,       --                    .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,           --                    .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,         --                    .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,         --                    .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,         --                    .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,        --                    .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready,        --                    .rready
			f2h_irq_p0               => hps_0_f2h_irq0_irq,                    --            f2h_irq0.irq
			f2h_irq_p1               => hps_0_f2h_irq1_irq                     --            f2h_irq1.irq
		);

	intr_capturer_0 : component intr_capturer
		generic map (
			NUM_INTR => 32
		)
		port map (
			clk          => pll_0_outclk0_clk,                                           --              clock.clk
			rst_n        => rst_controller_reset_out_reset_ports_inv,                    --         reset_sink.reset_n
			addr         => mm_interconnect_3_intr_capturer_0_avalon_slave_0_address(0), --     avalon_slave_0.address
			read         => mm_interconnect_3_intr_capturer_0_avalon_slave_0_read,       --                   .read
			rddata       => mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata,   --                   .readdata
			interrupt_in => intr_capturer_0_interrupt_receiver_irq                       -- interrupt_receiver.irq
		);

	lw_mm_bridge : component soc_system_lw_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 20,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => pll_0_outclk0_clk,                               --   clk.clk
			reset            => rst_controller_reset_out_reset,                  -- reset.reset
			s0_waitrequest   => mm_interconnect_2_lw_mm_bridge_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_interconnect_2_lw_mm_bridge_s0_readdata,      --      .readdata
			s0_readdatavalid => mm_interconnect_2_lw_mm_bridge_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_interconnect_2_lw_mm_bridge_s0_burstcount,    --      .burstcount
			s0_writedata     => mm_interconnect_2_lw_mm_bridge_s0_writedata,     --      .writedata
			s0_address       => mm_interconnect_2_lw_mm_bridge_s0_address,       --      .address
			s0_write         => mm_interconnect_2_lw_mm_bridge_s0_write,         --      .write
			s0_read          => mm_interconnect_2_lw_mm_bridge_s0_read,          --      .read
			s0_byteenable    => mm_interconnect_2_lw_mm_bridge_s0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_interconnect_2_lw_mm_bridge_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => lw_mm_bridge_m0_waitrequest,                     --    m0.waitrequest
			m0_readdata      => lw_mm_bridge_m0_readdata,                        --      .readdata
			m0_readdatavalid => lw_mm_bridge_m0_readdatavalid,                   --      .readdatavalid
			m0_burstcount    => lw_mm_bridge_m0_burstcount,                      --      .burstcount
			m0_writedata     => lw_mm_bridge_m0_writedata,                       --      .writedata
			m0_address       => lw_mm_bridge_m0_address,                         --      .address
			m0_write         => lw_mm_bridge_m0_write,                           --      .write
			m0_read          => lw_mm_bridge_m0_read,                            --      .read
			m0_byteenable    => lw_mm_bridge_m0_byteenable,                      --      .byteenable
			m0_debugaccess   => lw_mm_bridge_m0_debugaccess,                     --      .debugaccess
			s0_response      => open,                                            -- (terminated)
			m0_response      => "00"                                             -- (terminated)
		);

	pll_0 : component soc_system_pll_0
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,       -- outclk0.clk
			outclk_1 => pll_0_outclk1_clk,       -- outclk1.clk
			locked   => open                     -- (terminated)
		);

	sysid_qsys : component soc_system_sysid_qsys
		port map (
			clock    => pll_0_outclk0_clk,                                     --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_3_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_3_sysid_qsys_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			axi_bridge_for_acp_128_0_s0_awid                 => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awid,    --                axi_bridge_for_acp_128_0_s0.awid
			axi_bridge_for_acp_128_0_s0_awaddr               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awaddr,  --                                           .awaddr
			axi_bridge_for_acp_128_0_s0_awlen                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlen,   --                                           .awlen
			axi_bridge_for_acp_128_0_s0_awsize               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awsize,  --                                           .awsize
			axi_bridge_for_acp_128_0_s0_awburst              => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awburst, --                                           .awburst
			axi_bridge_for_acp_128_0_s0_awlock               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlock,  --                                           .awlock
			axi_bridge_for_acp_128_0_s0_awcache              => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awcache, --                                           .awcache
			axi_bridge_for_acp_128_0_s0_awprot               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awprot,  --                                           .awprot
			axi_bridge_for_acp_128_0_s0_awuser               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awuser,  --                                           .awuser
			axi_bridge_for_acp_128_0_s0_awvalid              => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awvalid, --                                           .awvalid
			axi_bridge_for_acp_128_0_s0_awready              => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awready, --                                           .awready
			axi_bridge_for_acp_128_0_s0_wid                  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wid,     --                                           .wid
			axi_bridge_for_acp_128_0_s0_wdata                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wdata,   --                                           .wdata
			axi_bridge_for_acp_128_0_s0_wstrb                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wstrb,   --                                           .wstrb
			axi_bridge_for_acp_128_0_s0_wlast                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wlast,   --                                           .wlast
			axi_bridge_for_acp_128_0_s0_wvalid               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wvalid,  --                                           .wvalid
			axi_bridge_for_acp_128_0_s0_wready               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wready,  --                                           .wready
			axi_bridge_for_acp_128_0_s0_bid                  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bid,     --                                           .bid
			axi_bridge_for_acp_128_0_s0_bresp                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bresp,   --                                           .bresp
			axi_bridge_for_acp_128_0_s0_bvalid               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bvalid,  --                                           .bvalid
			axi_bridge_for_acp_128_0_s0_bready               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bready,  --                                           .bready
			axi_bridge_for_acp_128_0_s0_arid                 => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arid,    --                                           .arid
			axi_bridge_for_acp_128_0_s0_araddr               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_araddr,  --                                           .araddr
			axi_bridge_for_acp_128_0_s0_arlen                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlen,   --                                           .arlen
			axi_bridge_for_acp_128_0_s0_arsize               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arsize,  --                                           .arsize
			axi_bridge_for_acp_128_0_s0_arburst              => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arburst, --                                           .arburst
			axi_bridge_for_acp_128_0_s0_arlock               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlock,  --                                           .arlock
			axi_bridge_for_acp_128_0_s0_arcache              => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arcache, --                                           .arcache
			axi_bridge_for_acp_128_0_s0_arprot               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arprot,  --                                           .arprot
			axi_bridge_for_acp_128_0_s0_aruser               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_aruser,  --                                           .aruser
			axi_bridge_for_acp_128_0_s0_arvalid              => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arvalid, --                                           .arvalid
			axi_bridge_for_acp_128_0_s0_arready              => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arready, --                                           .arready
			axi_bridge_for_acp_128_0_s0_rid                  => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rid,     --                                           .rid
			axi_bridge_for_acp_128_0_s0_rdata                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rdata,   --                                           .rdata
			axi_bridge_for_acp_128_0_s0_rresp                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rresp,   --                                           .rresp
			axi_bridge_for_acp_128_0_s0_rlast                => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rlast,   --                                           .rlast
			axi_bridge_for_acp_128_0_s0_rvalid               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rvalid,  --                                           .rvalid
			axi_bridge_for_acp_128_0_s0_rready               => mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rready,  --                                           .rready
			pll_0_outclk0_clk                                => pll_0_outclk0_clk,                                     --                              pll_0_outclk0.clk
			fft_ddr_bridge_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                        -- fft_ddr_bridge_reset_reset_bridge_in_reset.reset
			fft_ddr_bridge_expanded_master_address           => fft_ddr_bridge_expanded_master_address,                --             fft_ddr_bridge_expanded_master.address
			fft_ddr_bridge_expanded_master_waitrequest       => fft_ddr_bridge_expanded_master_waitrequest,            --                                           .waitrequest
			fft_ddr_bridge_expanded_master_burstcount        => fft_ddr_bridge_expanded_master_burstcount,             --                                           .burstcount
			fft_ddr_bridge_expanded_master_byteenable        => fft_ddr_bridge_expanded_master_byteenable,             --                                           .byteenable
			fft_ddr_bridge_expanded_master_read              => fft_ddr_bridge_expanded_master_read,                   --                                           .read
			fft_ddr_bridge_expanded_master_readdata          => fft_ddr_bridge_expanded_master_readdata,               --                                           .readdata
			fft_ddr_bridge_expanded_master_readdatavalid     => fft_ddr_bridge_expanded_master_readdatavalid,          --                                           .readdatavalid
			fft_ddr_bridge_expanded_master_write             => fft_ddr_bridge_expanded_master_write,                  --                                           .write
			fft_ddr_bridge_expanded_master_writedata         => fft_ddr_bridge_expanded_master_writedata               --                                           .writedata
		);

	mm_interconnect_1 : component soc_system_mm_interconnect_1
		port map (
			hps_0_h2f_axi_master_awid                                        => hps_0_h2f_axi_master_awid,                               --                                       hps_0_h2f_axi_master.awid
			hps_0_h2f_axi_master_awaddr                                      => hps_0_h2f_axi_master_awaddr,                             --                                                           .awaddr
			hps_0_h2f_axi_master_awlen                                       => hps_0_h2f_axi_master_awlen,                              --                                                           .awlen
			hps_0_h2f_axi_master_awsize                                      => hps_0_h2f_axi_master_awsize,                             --                                                           .awsize
			hps_0_h2f_axi_master_awburst                                     => hps_0_h2f_axi_master_awburst,                            --                                                           .awburst
			hps_0_h2f_axi_master_awlock                                      => hps_0_h2f_axi_master_awlock,                             --                                                           .awlock
			hps_0_h2f_axi_master_awcache                                     => hps_0_h2f_axi_master_awcache,                            --                                                           .awcache
			hps_0_h2f_axi_master_awprot                                      => hps_0_h2f_axi_master_awprot,                             --                                                           .awprot
			hps_0_h2f_axi_master_awvalid                                     => hps_0_h2f_axi_master_awvalid,                            --                                                           .awvalid
			hps_0_h2f_axi_master_awready                                     => hps_0_h2f_axi_master_awready,                            --                                                           .awready
			hps_0_h2f_axi_master_wid                                         => hps_0_h2f_axi_master_wid,                                --                                                           .wid
			hps_0_h2f_axi_master_wdata                                       => hps_0_h2f_axi_master_wdata,                              --                                                           .wdata
			hps_0_h2f_axi_master_wstrb                                       => hps_0_h2f_axi_master_wstrb,                              --                                                           .wstrb
			hps_0_h2f_axi_master_wlast                                       => hps_0_h2f_axi_master_wlast,                              --                                                           .wlast
			hps_0_h2f_axi_master_wvalid                                      => hps_0_h2f_axi_master_wvalid,                             --                                                           .wvalid
			hps_0_h2f_axi_master_wready                                      => hps_0_h2f_axi_master_wready,                             --                                                           .wready
			hps_0_h2f_axi_master_bid                                         => hps_0_h2f_axi_master_bid,                                --                                                           .bid
			hps_0_h2f_axi_master_bresp                                       => hps_0_h2f_axi_master_bresp,                              --                                                           .bresp
			hps_0_h2f_axi_master_bvalid                                      => hps_0_h2f_axi_master_bvalid,                             --                                                           .bvalid
			hps_0_h2f_axi_master_bready                                      => hps_0_h2f_axi_master_bready,                             --                                                           .bready
			hps_0_h2f_axi_master_arid                                        => hps_0_h2f_axi_master_arid,                               --                                                           .arid
			hps_0_h2f_axi_master_araddr                                      => hps_0_h2f_axi_master_araddr,                             --                                                           .araddr
			hps_0_h2f_axi_master_arlen                                       => hps_0_h2f_axi_master_arlen,                              --                                                           .arlen
			hps_0_h2f_axi_master_arsize                                      => hps_0_h2f_axi_master_arsize,                             --                                                           .arsize
			hps_0_h2f_axi_master_arburst                                     => hps_0_h2f_axi_master_arburst,                            --                                                           .arburst
			hps_0_h2f_axi_master_arlock                                      => hps_0_h2f_axi_master_arlock,                             --                                                           .arlock
			hps_0_h2f_axi_master_arcache                                     => hps_0_h2f_axi_master_arcache,                            --                                                           .arcache
			hps_0_h2f_axi_master_arprot                                      => hps_0_h2f_axi_master_arprot,                             --                                                           .arprot
			hps_0_h2f_axi_master_arvalid                                     => hps_0_h2f_axi_master_arvalid,                            --                                                           .arvalid
			hps_0_h2f_axi_master_arready                                     => hps_0_h2f_axi_master_arready,                            --                                                           .arready
			hps_0_h2f_axi_master_rid                                         => hps_0_h2f_axi_master_rid,                                --                                                           .rid
			hps_0_h2f_axi_master_rdata                                       => hps_0_h2f_axi_master_rdata,                              --                                                           .rdata
			hps_0_h2f_axi_master_rresp                                       => hps_0_h2f_axi_master_rresp,                              --                                                           .rresp
			hps_0_h2f_axi_master_rlast                                       => hps_0_h2f_axi_master_rlast,                              --                                                           .rlast
			hps_0_h2f_axi_master_rvalid                                      => hps_0_h2f_axi_master_rvalid,                             --                                                           .rvalid
			hps_0_h2f_axi_master_rready                                      => hps_0_h2f_axi_master_rready,                             --                                                           .rready
			pll_0_outclk0_clk                                                => pll_0_outclk0_clk,                                       --                                              pll_0_outclk0.clk
			FPGA_Slave_mm_bridge_reset_reset_bridge_in_reset_reset           => rst_controller_reset_out_reset,                          --           FPGA_Slave_mm_bridge_reset_reset_bridge_in_reset.reset
			hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                      -- hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			FPGA_Slave_mm_bridge_s0_address                                  => mm_interconnect_1_fpga_slave_mm_bridge_s0_address,       --                                    FPGA_Slave_mm_bridge_s0.address
			FPGA_Slave_mm_bridge_s0_write                                    => mm_interconnect_1_fpga_slave_mm_bridge_s0_write,         --                                                           .write
			FPGA_Slave_mm_bridge_s0_read                                     => mm_interconnect_1_fpga_slave_mm_bridge_s0_read,          --                                                           .read
			FPGA_Slave_mm_bridge_s0_readdata                                 => mm_interconnect_1_fpga_slave_mm_bridge_s0_readdata,      --                                                           .readdata
			FPGA_Slave_mm_bridge_s0_writedata                                => mm_interconnect_1_fpga_slave_mm_bridge_s0_writedata,     --                                                           .writedata
			FPGA_Slave_mm_bridge_s0_burstcount                               => mm_interconnect_1_fpga_slave_mm_bridge_s0_burstcount,    --                                                           .burstcount
			FPGA_Slave_mm_bridge_s0_byteenable                               => mm_interconnect_1_fpga_slave_mm_bridge_s0_byteenable,    --                                                           .byteenable
			FPGA_Slave_mm_bridge_s0_readdatavalid                            => mm_interconnect_1_fpga_slave_mm_bridge_s0_readdatavalid, --                                                           .readdatavalid
			FPGA_Slave_mm_bridge_s0_waitrequest                              => mm_interconnect_1_fpga_slave_mm_bridge_s0_waitrequest,   --                                                           .waitrequest
			FPGA_Slave_mm_bridge_s0_debugaccess                              => mm_interconnect_1_fpga_slave_mm_bridge_s0_debugaccess    --                                                           .debugaccess
		);

	mm_interconnect_2 : component soc_system_mm_interconnect_2
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                    --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                  --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                   --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                  --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                 --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                  --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                 --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                  --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                 --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                 --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                     --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                   --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                   --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                   --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                  --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                  --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                     --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                   --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                  --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                  --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                    --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                  --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                   --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                  --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                 --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                  --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                 --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                  --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                 --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                 --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                     --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                   --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                   --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                   --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                  --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                  --                                                              .rready
			pll_0_outclk0_clk                                                   => pll_0_outclk0_clk,                               --                                                 pll_0_outclk0.clk
			fpga_only_master_clk_reset_reset_bridge_in_reset_reset              => rst_controller_reset_out_reset,                  --              fpga_only_master_clk_reset_reset_bridge_in_reset.reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,              -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			lw_mm_bridge_reset_reset_bridge_in_reset_reset                      => rst_controller_reset_out_reset,                  --                      lw_mm_bridge_reset_reset_bridge_in_reset.reset
			fpga_only_master_master_address                                     => fpga_only_master_master_address,                 --                                       fpga_only_master_master.address
			fpga_only_master_master_waitrequest                                 => fpga_only_master_master_waitrequest,             --                                                              .waitrequest
			fpga_only_master_master_byteenable                                  => fpga_only_master_master_byteenable,              --                                                              .byteenable
			fpga_only_master_master_read                                        => fpga_only_master_master_read,                    --                                                              .read
			fpga_only_master_master_readdata                                    => fpga_only_master_master_readdata,                --                                                              .readdata
			fpga_only_master_master_readdatavalid                               => fpga_only_master_master_readdatavalid,           --                                                              .readdatavalid
			fpga_only_master_master_write                                       => fpga_only_master_master_write,                   --                                                              .write
			fpga_only_master_master_writedata                                   => fpga_only_master_master_writedata,               --                                                              .writedata
			lw_mm_bridge_s0_address                                             => mm_interconnect_2_lw_mm_bridge_s0_address,       --                                               lw_mm_bridge_s0.address
			lw_mm_bridge_s0_write                                               => mm_interconnect_2_lw_mm_bridge_s0_write,         --                                                              .write
			lw_mm_bridge_s0_read                                                => mm_interconnect_2_lw_mm_bridge_s0_read,          --                                                              .read
			lw_mm_bridge_s0_readdata                                            => mm_interconnect_2_lw_mm_bridge_s0_readdata,      --                                                              .readdata
			lw_mm_bridge_s0_writedata                                           => mm_interconnect_2_lw_mm_bridge_s0_writedata,     --                                                              .writedata
			lw_mm_bridge_s0_burstcount                                          => mm_interconnect_2_lw_mm_bridge_s0_burstcount,    --                                                              .burstcount
			lw_mm_bridge_s0_byteenable                                          => mm_interconnect_2_lw_mm_bridge_s0_byteenable,    --                                                              .byteenable
			lw_mm_bridge_s0_readdatavalid                                       => mm_interconnect_2_lw_mm_bridge_s0_readdatavalid, --                                                              .readdatavalid
			lw_mm_bridge_s0_waitrequest                                         => mm_interconnect_2_lw_mm_bridge_s0_waitrequest,   --                                                              .waitrequest
			lw_mm_bridge_s0_debugaccess                                         => mm_interconnect_2_lw_mm_bridge_s0_debugaccess    --                                                              .debugaccess
		);

	mm_interconnect_3 : component soc_system_mm_interconnect_3
		port map (
			pll_0_outclk0_clk                              => pll_0_outclk0_clk,                                         --                            pll_0_outclk0.clk
			KBandIPsub_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                            --   KBandIPsub_reset_reset_bridge_in_reset.reset
			lw_mm_bridge_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- lw_mm_bridge_reset_reset_bridge_in_reset.reset
			lw_mm_bridge_m0_address                        => lw_mm_bridge_m0_address,                                   --                          lw_mm_bridge_m0.address
			lw_mm_bridge_m0_waitrequest                    => lw_mm_bridge_m0_waitrequest,                               --                                         .waitrequest
			lw_mm_bridge_m0_burstcount                     => lw_mm_bridge_m0_burstcount,                                --                                         .burstcount
			lw_mm_bridge_m0_byteenable                     => lw_mm_bridge_m0_byteenable,                                --                                         .byteenable
			lw_mm_bridge_m0_read                           => lw_mm_bridge_m0_read,                                      --                                         .read
			lw_mm_bridge_m0_readdata                       => lw_mm_bridge_m0_readdata,                                  --                                         .readdata
			lw_mm_bridge_m0_readdatavalid                  => lw_mm_bridge_m0_readdatavalid,                             --                                         .readdatavalid
			lw_mm_bridge_m0_write                          => lw_mm_bridge_m0_write,                                     --                                         .write
			lw_mm_bridge_m0_writedata                      => lw_mm_bridge_m0_writedata,                                 --                                         .writedata
			lw_mm_bridge_m0_debugaccess                    => lw_mm_bridge_m0_debugaccess,                               --                                         .debugaccess
			intr_capturer_0_avalon_slave_0_address         => mm_interconnect_3_intr_capturer_0_avalon_slave_0_address,  --           intr_capturer_0_avalon_slave_0.address
			intr_capturer_0_avalon_slave_0_read            => mm_interconnect_3_intr_capturer_0_avalon_slave_0_read,     --                                         .read
			intr_capturer_0_avalon_slave_0_readdata        => mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata, --                                         .readdata
			KBandIPsub_slw_address                         => mm_interconnect_3_kbandipsub_slw_address,                  --                           KBandIPsub_slw.address
			KBandIPsub_slw_write                           => mm_interconnect_3_kbandipsub_slw_write,                    --                                         .write
			KBandIPsub_slw_read                            => mm_interconnect_3_kbandipsub_slw_read,                     --                                         .read
			KBandIPsub_slw_readdata                        => mm_interconnect_3_kbandipsub_slw_readdata,                 --                                         .readdata
			KBandIPsub_slw_writedata                       => mm_interconnect_3_kbandipsub_slw_writedata,                --                                         .writedata
			KBandIPsub_slw_burstcount                      => mm_interconnect_3_kbandipsub_slw_burstcount,               --                                         .burstcount
			KBandIPsub_slw_byteenable                      => mm_interconnect_3_kbandipsub_slw_byteenable,               --                                         .byteenable
			KBandIPsub_slw_readdatavalid                   => mm_interconnect_3_kbandipsub_slw_readdatavalid,            --                                         .readdatavalid
			KBandIPsub_slw_waitrequest                     => mm_interconnect_3_kbandipsub_slw_waitrequest,              --                                         .waitrequest
			KBandIPsub_slw_debugaccess                     => mm_interconnect_3_kbandipsub_slw_debugaccess,              --                                         .debugaccess
			sysid_qsys_control_slave_address               => mm_interconnect_3_sysid_qsys_control_slave_address,        --                 sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata              => mm_interconnect_3_sysid_qsys_control_slave_readdata        --                                         .readdata
		);

	mm_interconnect_6 : component soc_system_mm_interconnect_6
		port map (
			pll_0_outclk0_clk                                => pll_0_outclk0_clk,                                             --                              pll_0_outclk0.clk
			fft_ddr_bridge_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                -- fft_ddr_bridge_reset_reset_bridge_in_reset.reset
			KBandIPsub_reset_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,                                --     KBandIPsub_reset_reset_bridge_in_reset.reset
			KBandIPsub_m0_address                            => kbandipsub_m0_address,                                         --                              KBandIPsub_m0.address
			KBandIPsub_m0_waitrequest                        => kbandipsub_m0_waitrequest,                                     --                                           .waitrequest
			KBandIPsub_m0_burstcount                         => kbandipsub_m0_burstcount,                                      --                                           .burstcount
			KBandIPsub_m0_byteenable                         => kbandipsub_m0_byteenable,                                      --                                           .byteenable
			KBandIPsub_m0_read                               => kbandipsub_m0_read,                                            --                                           .read
			KBandIPsub_m0_readdata                           => kbandipsub_m0_readdata,                                        --                                           .readdata
			KBandIPsub_m0_readdatavalid                      => kbandipsub_m0_readdatavalid,                                   --                                           .readdatavalid
			KBandIPsub_m0_write                              => kbandipsub_m0_write,                                           --                                           .write
			KBandIPsub_m0_writedata                          => kbandipsub_m0_writedata,                                       --                                           .writedata
			KBandIPsub_m0_debugaccess                        => kbandipsub_m0_debugaccess,                                     --                                           .debugaccess
			fft_ddr_bridge_windowed_slave_address            => mm_interconnect_6_fft_ddr_bridge_windowed_slave_address,       --              fft_ddr_bridge_windowed_slave.address
			fft_ddr_bridge_windowed_slave_write              => mm_interconnect_6_fft_ddr_bridge_windowed_slave_write,         --                                           .write
			fft_ddr_bridge_windowed_slave_read               => mm_interconnect_6_fft_ddr_bridge_windowed_slave_read,          --                                           .read
			fft_ddr_bridge_windowed_slave_readdata           => mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdata,      --                                           .readdata
			fft_ddr_bridge_windowed_slave_writedata          => mm_interconnect_6_fft_ddr_bridge_windowed_slave_writedata,     --                                           .writedata
			fft_ddr_bridge_windowed_slave_burstcount         => mm_interconnect_6_fft_ddr_bridge_windowed_slave_burstcount,    --                                           .burstcount
			fft_ddr_bridge_windowed_slave_byteenable         => mm_interconnect_6_fft_ddr_bridge_windowed_slave_byteenable,    --                                           .byteenable
			fft_ddr_bridge_windowed_slave_readdatavalid      => mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdatavalid, --                                           .readdatavalid
			fft_ddr_bridge_windowed_slave_waitrequest        => mm_interconnect_6_fft_ddr_bridge_windowed_slave_waitrequest    --                                           .waitrequest
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq, -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq, -- receiver2.irq
			sender_irq    => hps_0_f2h_irq0_irq        --    sender.irq
		);

	irq_mapper_001 : component soc_system_irq_mapper_001
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq1_irq  --    sender.irq
		);

	irq_mapper_002 : component soc_system_irq_mapper
		port map (
			clk           => pll_0_outclk0_clk,                      --       clk.clk
			reset         => rst_controller_reset_out_reset,         -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,               -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,               -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,               -- receiver2.irq
			sender_irq    => intr_capturer_0_interrupt_receiver_irq  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => pll_0_outclk0_clk,              --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_n_ports_inv,  -- reset_in0.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	hps_0_h2f_reset_reset_n_ports_inv <= not hps_0_h2f_reset_reset;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_n <= hps_0_h2f_reset_reset;

end architecture rtl; -- of soc_system
